
module fpMultiplier_DW01_add_2 ( A, B, CI, SUM, CO );
  input [45:0] A;
  input [45:0] B;
  output [45:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113;
  assign SUM[22] = A[22];
  assign SUM[21] = A[21];

  AND2_X1 U2 ( .A1(n2), .A2(n113), .ZN(SUM[23]) );
  OR2_X1 U3 ( .A1(B[23]), .A2(A[23]), .ZN(n2) );
  INV_X1 U4 ( .A(n34), .ZN(n8) );
  INV_X1 U5 ( .A(n104), .ZN(n25) );
  INV_X1 U6 ( .A(n96), .ZN(n23) );
  INV_X1 U7 ( .A(n88), .ZN(n21) );
  INV_X1 U8 ( .A(n80), .ZN(n19) );
  INV_X1 U9 ( .A(n64), .ZN(n15) );
  INV_X1 U10 ( .A(n56), .ZN(n13) );
  INV_X1 U11 ( .A(n48), .ZN(n11) );
  INV_X1 U12 ( .A(n40), .ZN(n9) );
  INV_X1 U13 ( .A(n32), .ZN(n7) );
  INV_X1 U14 ( .A(n72), .ZN(n17) );
  INV_X1 U15 ( .A(n42), .ZN(n10) );
  INV_X1 U16 ( .A(n106), .ZN(n26) );
  INV_X1 U17 ( .A(n98), .ZN(n24) );
  INV_X1 U18 ( .A(n90), .ZN(n22) );
  INV_X1 U19 ( .A(n82), .ZN(n20) );
  INV_X1 U20 ( .A(n74), .ZN(n18) );
  INV_X1 U21 ( .A(n58), .ZN(n14) );
  INV_X1 U22 ( .A(n50), .ZN(n12) );
  INV_X1 U23 ( .A(n66), .ZN(n16) );
  INV_X1 U24 ( .A(n111), .ZN(n27) );
  NAND2_X1 U25 ( .A1(n5), .A2(n6), .ZN(SUM[45]) );
  NAND2_X1 U26 ( .A1(B[45]), .A2(n29), .ZN(n5) );
  NAND2_X1 U27 ( .A1(n3), .A2(n4), .ZN(n6) );
  INV_X1 U28 ( .A(B[45]), .ZN(n3) );
  INV_X1 U29 ( .A(n29), .ZN(n4) );
  INV_X1 U30 ( .A(n113), .ZN(n28) );
  AOI21_X1 U31 ( .B1(n30), .B2(n7), .A(n31), .ZN(n29) );
  XOR2_X1 U32 ( .A(n30), .B(n33), .Z(SUM[44]) );
  NOR2_X1 U33 ( .A1(n31), .A2(n32), .ZN(n33) );
  NOR2_X1 U34 ( .A1(B[44]), .A2(A[44]), .ZN(n32) );
  AND2_X1 U35 ( .A1(B[44]), .A2(A[44]), .ZN(n31) );
  OAI21_X1 U36 ( .B1(n34), .B2(n35), .A(n36), .ZN(n30) );
  XOR2_X1 U37 ( .A(n37), .B(n35), .Z(SUM[43]) );
  AOI21_X1 U38 ( .B1(n9), .B2(n38), .A(n39), .ZN(n35) );
  NAND2_X1 U39 ( .A1(n8), .A2(n36), .ZN(n37) );
  NAND2_X1 U40 ( .A1(B[43]), .A2(A[43]), .ZN(n36) );
  NOR2_X1 U41 ( .A1(B[43]), .A2(A[43]), .ZN(n34) );
  XOR2_X1 U42 ( .A(n38), .B(n41), .Z(SUM[42]) );
  NOR2_X1 U43 ( .A1(n39), .A2(n40), .ZN(n41) );
  NOR2_X1 U44 ( .A1(B[42]), .A2(A[42]), .ZN(n40) );
  AND2_X1 U45 ( .A1(B[42]), .A2(A[42]), .ZN(n39) );
  OAI21_X1 U46 ( .B1(n42), .B2(n43), .A(n44), .ZN(n38) );
  XOR2_X1 U47 ( .A(n45), .B(n43), .Z(SUM[41]) );
  AOI21_X1 U48 ( .B1(n11), .B2(n46), .A(n47), .ZN(n43) );
  NAND2_X1 U49 ( .A1(n10), .A2(n44), .ZN(n45) );
  NAND2_X1 U50 ( .A1(B[41]), .A2(A[41]), .ZN(n44) );
  NOR2_X1 U51 ( .A1(B[41]), .A2(A[41]), .ZN(n42) );
  XOR2_X1 U52 ( .A(n46), .B(n49), .Z(SUM[40]) );
  NOR2_X1 U53 ( .A1(n47), .A2(n48), .ZN(n49) );
  NOR2_X1 U54 ( .A1(B[40]), .A2(A[40]), .ZN(n48) );
  AND2_X1 U55 ( .A1(B[40]), .A2(A[40]), .ZN(n47) );
  OAI21_X1 U56 ( .B1(n50), .B2(n51), .A(n52), .ZN(n46) );
  XOR2_X1 U57 ( .A(n53), .B(n51), .Z(SUM[39]) );
  AOI21_X1 U58 ( .B1(n13), .B2(n54), .A(n55), .ZN(n51) );
  NAND2_X1 U59 ( .A1(n12), .A2(n52), .ZN(n53) );
  NAND2_X1 U60 ( .A1(B[39]), .A2(A[39]), .ZN(n52) );
  NOR2_X1 U61 ( .A1(B[39]), .A2(A[39]), .ZN(n50) );
  XOR2_X1 U62 ( .A(n54), .B(n57), .Z(SUM[38]) );
  NOR2_X1 U63 ( .A1(n55), .A2(n56), .ZN(n57) );
  NOR2_X1 U64 ( .A1(B[38]), .A2(A[38]), .ZN(n56) );
  AND2_X1 U65 ( .A1(B[38]), .A2(A[38]), .ZN(n55) );
  OAI21_X1 U66 ( .B1(n58), .B2(n59), .A(n60), .ZN(n54) );
  XOR2_X1 U67 ( .A(n61), .B(n59), .Z(SUM[37]) );
  AOI21_X1 U68 ( .B1(n15), .B2(n62), .A(n63), .ZN(n59) );
  NAND2_X1 U69 ( .A1(n14), .A2(n60), .ZN(n61) );
  NAND2_X1 U70 ( .A1(B[37]), .A2(A[37]), .ZN(n60) );
  NOR2_X1 U71 ( .A1(B[37]), .A2(A[37]), .ZN(n58) );
  XOR2_X1 U72 ( .A(n62), .B(n65), .Z(SUM[36]) );
  NOR2_X1 U73 ( .A1(n63), .A2(n64), .ZN(n65) );
  NOR2_X1 U74 ( .A1(B[36]), .A2(A[36]), .ZN(n64) );
  AND2_X1 U75 ( .A1(B[36]), .A2(A[36]), .ZN(n63) );
  OAI21_X1 U76 ( .B1(n66), .B2(n67), .A(n68), .ZN(n62) );
  XOR2_X1 U77 ( .A(n69), .B(n67), .Z(SUM[35]) );
  AOI21_X1 U78 ( .B1(n17), .B2(n70), .A(n71), .ZN(n67) );
  NAND2_X1 U79 ( .A1(n16), .A2(n68), .ZN(n69) );
  NAND2_X1 U80 ( .A1(B[35]), .A2(A[35]), .ZN(n68) );
  NOR2_X1 U81 ( .A1(B[35]), .A2(A[35]), .ZN(n66) );
  XOR2_X1 U82 ( .A(n70), .B(n73), .Z(SUM[34]) );
  NOR2_X1 U83 ( .A1(n71), .A2(n72), .ZN(n73) );
  NOR2_X1 U84 ( .A1(B[34]), .A2(A[34]), .ZN(n72) );
  AND2_X1 U85 ( .A1(B[34]), .A2(A[34]), .ZN(n71) );
  OAI21_X1 U86 ( .B1(n74), .B2(n75), .A(n76), .ZN(n70) );
  XOR2_X1 U87 ( .A(n77), .B(n75), .Z(SUM[33]) );
  AOI21_X1 U88 ( .B1(n19), .B2(n78), .A(n79), .ZN(n75) );
  NAND2_X1 U89 ( .A1(n18), .A2(n76), .ZN(n77) );
  NAND2_X1 U90 ( .A1(B[33]), .A2(A[33]), .ZN(n76) );
  NOR2_X1 U91 ( .A1(B[33]), .A2(A[33]), .ZN(n74) );
  XOR2_X1 U92 ( .A(n78), .B(n81), .Z(SUM[32]) );
  NOR2_X1 U93 ( .A1(n79), .A2(n80), .ZN(n81) );
  NOR2_X1 U94 ( .A1(B[32]), .A2(A[32]), .ZN(n80) );
  AND2_X1 U95 ( .A1(B[32]), .A2(A[32]), .ZN(n79) );
  OAI21_X1 U96 ( .B1(n82), .B2(n83), .A(n84), .ZN(n78) );
  XOR2_X1 U97 ( .A(n85), .B(n83), .Z(SUM[31]) );
  AOI21_X1 U98 ( .B1(n21), .B2(n86), .A(n87), .ZN(n83) );
  NAND2_X1 U99 ( .A1(n20), .A2(n84), .ZN(n85) );
  NAND2_X1 U100 ( .A1(B[31]), .A2(A[31]), .ZN(n84) );
  NOR2_X1 U101 ( .A1(B[31]), .A2(A[31]), .ZN(n82) );
  XOR2_X1 U102 ( .A(n86), .B(n89), .Z(SUM[30]) );
  NOR2_X1 U103 ( .A1(n87), .A2(n88), .ZN(n89) );
  NOR2_X1 U104 ( .A1(B[30]), .A2(A[30]), .ZN(n88) );
  AND2_X1 U105 ( .A1(B[30]), .A2(A[30]), .ZN(n87) );
  OAI21_X1 U106 ( .B1(n90), .B2(n91), .A(n92), .ZN(n86) );
  XOR2_X1 U107 ( .A(n93), .B(n91), .Z(SUM[29]) );
  AOI21_X1 U108 ( .B1(n23), .B2(n94), .A(n95), .ZN(n91) );
  NAND2_X1 U109 ( .A1(n22), .A2(n92), .ZN(n93) );
  NAND2_X1 U110 ( .A1(B[29]), .A2(A[29]), .ZN(n92) );
  NOR2_X1 U111 ( .A1(B[29]), .A2(A[29]), .ZN(n90) );
  XOR2_X1 U112 ( .A(n94), .B(n97), .Z(SUM[28]) );
  NOR2_X1 U113 ( .A1(n95), .A2(n96), .ZN(n97) );
  NOR2_X1 U114 ( .A1(B[28]), .A2(A[28]), .ZN(n96) );
  AND2_X1 U115 ( .A1(B[28]), .A2(A[28]), .ZN(n95) );
  OAI21_X1 U116 ( .B1(n98), .B2(n99), .A(n100), .ZN(n94) );
  XOR2_X1 U117 ( .A(n101), .B(n99), .Z(SUM[27]) );
  AOI21_X1 U118 ( .B1(n102), .B2(n25), .A(n103), .ZN(n99) );
  NAND2_X1 U119 ( .A1(n24), .A2(n100), .ZN(n101) );
  NAND2_X1 U120 ( .A1(B[27]), .A2(A[27]), .ZN(n100) );
  NOR2_X1 U121 ( .A1(B[27]), .A2(A[27]), .ZN(n98) );
  XOR2_X1 U122 ( .A(n102), .B(n105), .Z(SUM[26]) );
  NOR2_X1 U123 ( .A1(n103), .A2(n104), .ZN(n105) );
  NOR2_X1 U124 ( .A1(B[26]), .A2(A[26]), .ZN(n104) );
  AND2_X1 U125 ( .A1(B[26]), .A2(A[26]), .ZN(n103) );
  OAI21_X1 U126 ( .B1(n106), .B2(n107), .A(n108), .ZN(n102) );
  XOR2_X1 U127 ( .A(n109), .B(n107), .Z(SUM[25]) );
  AOI21_X1 U128 ( .B1(n27), .B2(n28), .A(n110), .ZN(n107) );
  NAND2_X1 U129 ( .A1(n26), .A2(n108), .ZN(n109) );
  NAND2_X1 U130 ( .A1(B[25]), .A2(A[25]), .ZN(n108) );
  NOR2_X1 U131 ( .A1(B[25]), .A2(A[25]), .ZN(n106) );
  XOR2_X1 U132 ( .A(n28), .B(n112), .Z(SUM[24]) );
  NOR2_X1 U133 ( .A1(n110), .A2(n111), .ZN(n112) );
  NOR2_X1 U134 ( .A1(B[24]), .A2(A[24]), .ZN(n111) );
  AND2_X1 U135 ( .A1(B[24]), .A2(A[24]), .ZN(n110) );
  NAND2_X1 U136 ( .A1(B[23]), .A2(A[23]), .ZN(n113) );
endmodule


module fpMultiplier_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [23:0] A;
  input [23:0] B;
  output [47:0] PRODUCT;
  input TC;
  wire   ab_23__23_, ab_23__22_, ab_23__21_, ab_23__20_, ab_23__19_,
         ab_23__18_, ab_23__17_, ab_23__16_, ab_23__15_, ab_23__14_,
         ab_23__13_, ab_23__12_, ab_23__11_, ab_23__10_, ab_23__9_, ab_23__8_,
         ab_23__7_, ab_23__6_, ab_23__5_, ab_23__4_, ab_23__3_, ab_23__2_,
         ab_23__1_, ab_23__0_, ab_22__23_, ab_22__22_, ab_22__21_, ab_22__20_,
         ab_22__19_, ab_22__18_, ab_22__17_, ab_22__16_, ab_22__15_,
         ab_22__14_, ab_22__13_, ab_22__12_, ab_22__11_, ab_22__10_, ab_22__9_,
         ab_22__8_, ab_22__7_, ab_22__6_, ab_22__5_, ab_22__4_, ab_22__3_,
         ab_22__2_, ab_22__1_, ab_22__0_, ab_21__23_, ab_21__22_, ab_21__21_,
         ab_21__20_, ab_21__19_, ab_21__18_, ab_21__17_, ab_21__16_,
         ab_21__15_, ab_21__14_, ab_21__13_, ab_21__12_, ab_21__11_,
         ab_21__10_, ab_21__9_, ab_21__8_, ab_21__7_, ab_21__6_, ab_21__5_,
         ab_21__4_, ab_21__3_, ab_21__2_, ab_21__1_, ab_21__0_, ab_20__23_,
         ab_20__22_, ab_20__21_, ab_20__20_, ab_20__19_, ab_20__18_,
         ab_20__17_, ab_20__16_, ab_20__15_, ab_20__14_, ab_20__13_,
         ab_20__12_, ab_20__11_, ab_20__10_, ab_20__9_, ab_20__8_, ab_20__7_,
         ab_20__6_, ab_20__5_, ab_20__4_, ab_20__3_, ab_20__2_, ab_20__1_,
         ab_20__0_, ab_19__23_, ab_19__22_, ab_19__21_, ab_19__20_, ab_19__19_,
         ab_19__18_, ab_19__17_, ab_19__16_, ab_19__15_, ab_19__14_,
         ab_19__13_, ab_19__12_, ab_19__11_, ab_19__10_, ab_19__9_, ab_19__8_,
         ab_19__7_, ab_19__6_, ab_19__5_, ab_19__4_, ab_19__3_, ab_19__2_,
         ab_19__1_, ab_19__0_, ab_18__23_, ab_18__22_, ab_18__21_, ab_18__20_,
         ab_18__19_, ab_18__18_, ab_18__17_, ab_18__16_, ab_18__15_,
         ab_18__14_, ab_18__13_, ab_18__12_, ab_18__11_, ab_18__10_, ab_18__9_,
         ab_18__8_, ab_18__7_, ab_18__6_, ab_18__5_, ab_18__4_, ab_18__3_,
         ab_18__2_, ab_18__1_, ab_18__0_, ab_17__23_, ab_17__22_, ab_17__21_,
         ab_17__20_, ab_17__19_, ab_17__18_, ab_17__17_, ab_17__16_,
         ab_17__15_, ab_17__14_, ab_17__13_, ab_17__12_, ab_17__11_,
         ab_17__10_, ab_17__9_, ab_17__8_, ab_17__7_, ab_17__6_, ab_17__5_,
         ab_17__4_, ab_17__3_, ab_17__2_, ab_17__1_, ab_17__0_, ab_16__23_,
         ab_16__22_, ab_16__21_, ab_16__20_, ab_16__19_, ab_16__18_,
         ab_16__17_, ab_16__16_, ab_16__15_, ab_16__14_, ab_16__13_,
         ab_16__12_, ab_16__11_, ab_16__10_, ab_16__9_, ab_16__8_, ab_16__7_,
         ab_16__6_, ab_16__5_, ab_16__4_, ab_16__3_, ab_16__2_, ab_16__1_,
         ab_16__0_, ab_15__23_, ab_15__22_, ab_15__21_, ab_15__20_, ab_15__19_,
         ab_15__18_, ab_15__17_, ab_15__16_, ab_15__15_, ab_15__14_,
         ab_15__13_, ab_15__12_, ab_15__11_, ab_15__10_, ab_15__9_, ab_15__8_,
         ab_15__7_, ab_15__6_, ab_15__5_, ab_15__4_, ab_15__3_, ab_15__2_,
         ab_15__1_, ab_15__0_, ab_14__23_, ab_14__22_, ab_14__21_, ab_14__20_,
         ab_14__19_, ab_14__18_, ab_14__17_, ab_14__16_, ab_14__15_,
         ab_14__14_, ab_14__13_, ab_14__12_, ab_14__11_, ab_14__10_, ab_14__9_,
         ab_14__8_, ab_14__7_, ab_14__6_, ab_14__5_, ab_14__4_, ab_14__3_,
         ab_14__2_, ab_14__1_, ab_14__0_, ab_13__23_, ab_13__22_, ab_13__21_,
         ab_13__20_, ab_13__19_, ab_13__18_, ab_13__17_, ab_13__16_,
         ab_13__15_, ab_13__14_, ab_13__13_, ab_13__12_, ab_13__11_,
         ab_13__10_, ab_13__9_, ab_13__8_, ab_13__7_, ab_13__6_, ab_13__5_,
         ab_13__4_, ab_13__3_, ab_13__2_, ab_13__1_, ab_13__0_, ab_12__23_,
         ab_12__22_, ab_12__21_, ab_12__20_, ab_12__19_, ab_12__18_,
         ab_12__17_, ab_12__16_, ab_12__15_, ab_12__14_, ab_12__13_,
         ab_12__12_, ab_12__11_, ab_12__10_, ab_12__9_, ab_12__8_, ab_12__7_,
         ab_12__6_, ab_12__5_, ab_12__4_, ab_12__3_, ab_12__2_, ab_12__1_,
         ab_12__0_, ab_11__23_, ab_11__22_, ab_11__21_, ab_11__20_, ab_11__19_,
         ab_11__18_, ab_11__17_, ab_11__16_, ab_11__15_, ab_11__14_,
         ab_11__13_, ab_11__12_, ab_11__11_, ab_11__10_, ab_11__9_, ab_11__8_,
         ab_11__7_, ab_11__6_, ab_11__5_, ab_11__4_, ab_11__3_, ab_11__2_,
         ab_11__1_, ab_11__0_, ab_10__23_, ab_10__22_, ab_10__21_, ab_10__20_,
         ab_10__19_, ab_10__18_, ab_10__17_, ab_10__16_, ab_10__15_,
         ab_10__14_, ab_10__13_, ab_10__12_, ab_10__11_, ab_10__10_, ab_10__9_,
         ab_10__8_, ab_10__7_, ab_10__6_, ab_10__5_, ab_10__4_, ab_10__3_,
         ab_10__2_, ab_10__1_, ab_10__0_, ab_9__23_, ab_9__22_, ab_9__21_,
         ab_9__20_, ab_9__19_, ab_9__18_, ab_9__17_, ab_9__16_, ab_9__15_,
         ab_9__14_, ab_9__13_, ab_9__12_, ab_9__11_, ab_9__10_, ab_9__9_,
         ab_9__8_, ab_9__7_, ab_9__6_, ab_9__5_, ab_9__4_, ab_9__3_, ab_9__2_,
         ab_9__1_, ab_9__0_, ab_8__23_, ab_8__22_, ab_8__21_, ab_8__20_,
         ab_8__19_, ab_8__18_, ab_8__17_, ab_8__16_, ab_8__15_, ab_8__14_,
         ab_8__13_, ab_8__12_, ab_8__11_, ab_8__10_, ab_8__9_, ab_8__8_,
         ab_8__7_, ab_8__6_, ab_8__5_, ab_8__4_, ab_8__3_, ab_8__2_, ab_8__1_,
         ab_8__0_, ab_7__23_, ab_7__22_, ab_7__21_, ab_7__20_, ab_7__19_,
         ab_7__18_, ab_7__17_, ab_7__16_, ab_7__15_, ab_7__14_, ab_7__13_,
         ab_7__12_, ab_7__11_, ab_7__10_, ab_7__9_, ab_7__8_, ab_7__7_,
         ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_, ab_7__0_,
         ab_6__23_, ab_6__22_, ab_6__21_, ab_6__20_, ab_6__19_, ab_6__18_,
         ab_6__17_, ab_6__16_, ab_6__15_, ab_6__14_, ab_6__13_, ab_6__12_,
         ab_6__11_, ab_6__10_, ab_6__9_, ab_6__8_, ab_6__7_, ab_6__6_,
         ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_, ab_6__1_, ab_6__0_, ab_5__23_,
         ab_5__22_, ab_5__21_, ab_5__20_, ab_5__19_, ab_5__18_, ab_5__17_,
         ab_5__16_, ab_5__15_, ab_5__14_, ab_5__13_, ab_5__12_, ab_5__11_,
         ab_5__10_, ab_5__9_, ab_5__8_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_,
         ab_5__3_, ab_5__2_, ab_5__1_, ab_5__0_, ab_4__23_, ab_4__22_,
         ab_4__21_, ab_4__20_, ab_4__19_, ab_4__18_, ab_4__17_, ab_4__16_,
         ab_4__15_, ab_4__14_, ab_4__13_, ab_4__12_, ab_4__11_, ab_4__10_,
         ab_4__9_, ab_4__8_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_, ab_4__3_,
         ab_4__2_, ab_4__1_, ab_4__0_, ab_3__23_, ab_3__22_, ab_3__21_,
         ab_3__20_, ab_3__19_, ab_3__18_, ab_3__17_, ab_3__16_, ab_3__15_,
         ab_3__14_, ab_3__13_, ab_3__12_, ab_3__11_, ab_3__10_, ab_3__9_,
         ab_3__8_, ab_3__7_, ab_3__6_, ab_3__5_, ab_3__4_, ab_3__3_, ab_3__2_,
         ab_3__1_, ab_3__0_, ab_2__23_, ab_2__22_, ab_2__21_, ab_2__20_,
         ab_2__19_, ab_2__18_, ab_2__17_, ab_2__16_, ab_2__15_, ab_2__14_,
         ab_2__13_, ab_2__12_, ab_2__11_, ab_2__10_, ab_2__9_, ab_2__8_,
         ab_2__7_, ab_2__6_, ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_,
         ab_2__0_, ab_1__23_, ab_1__22_, ab_1__21_, ab_1__20_, ab_1__19_,
         ab_1__18_, ab_1__17_, ab_1__16_, ab_1__15_, ab_1__14_, ab_1__13_,
         ab_1__12_, ab_1__11_, ab_1__10_, ab_1__9_, ab_1__8_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_0__23_,
         ab_0__22_, ab_0__21_, ab_0__20_, ab_0__19_, ab_0__18_, ab_0__17_,
         ab_0__16_, ab_0__15_, ab_0__14_, ab_0__13_, ab_0__12_, ab_0__11_,
         ab_0__10_, ab_0__9_, ab_0__8_, ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_,
         ab_0__3_, ab_0__2_, CARRYB_23__22_, CARRYB_23__21_, CARRYB_23__20_,
         CARRYB_23__19_, CARRYB_23__18_, CARRYB_23__17_, CARRYB_23__16_,
         CARRYB_23__15_, CARRYB_23__14_, CARRYB_23__13_, CARRYB_23__12_,
         CARRYB_23__11_, CARRYB_23__10_, CARRYB_23__9_, CARRYB_23__8_,
         CARRYB_23__7_, CARRYB_23__6_, CARRYB_23__5_, CARRYB_23__4_,
         CARRYB_23__3_, CARRYB_23__2_, CARRYB_23__1_, CARRYB_23__0_,
         CARRYB_22__22_, CARRYB_22__21_, CARRYB_22__20_, CARRYB_22__19_,
         CARRYB_22__18_, CARRYB_22__17_, CARRYB_22__16_, CARRYB_22__15_,
         CARRYB_22__14_, CARRYB_22__13_, CARRYB_22__12_, CARRYB_22__11_,
         CARRYB_22__10_, CARRYB_22__9_, CARRYB_22__8_, CARRYB_22__7_,
         CARRYB_22__6_, CARRYB_22__5_, CARRYB_22__4_, CARRYB_22__3_,
         CARRYB_22__2_, CARRYB_22__1_, CARRYB_22__0_, CARRYB_21__22_,
         CARRYB_21__21_, CARRYB_21__20_, CARRYB_21__19_, CARRYB_21__18_,
         CARRYB_21__17_, CARRYB_21__16_, CARRYB_21__15_, CARRYB_21__14_,
         CARRYB_21__13_, CARRYB_21__12_, CARRYB_21__11_, CARRYB_21__10_,
         CARRYB_21__9_, CARRYB_21__8_, CARRYB_21__7_, CARRYB_21__6_,
         CARRYB_21__5_, CARRYB_21__4_, CARRYB_21__3_, CARRYB_21__2_,
         CARRYB_21__1_, CARRYB_21__0_, CARRYB_20__22_, CARRYB_20__21_,
         CARRYB_20__20_, CARRYB_20__19_, CARRYB_20__18_, CARRYB_20__17_,
         CARRYB_20__16_, CARRYB_20__15_, CARRYB_20__14_, CARRYB_20__13_,
         CARRYB_20__12_, CARRYB_20__11_, CARRYB_20__10_, CARRYB_20__9_,
         CARRYB_20__8_, CARRYB_20__7_, CARRYB_20__6_, CARRYB_20__5_,
         CARRYB_20__4_, CARRYB_20__3_, CARRYB_20__2_, CARRYB_20__1_,
         CARRYB_20__0_, CARRYB_19__22_, CARRYB_19__21_, CARRYB_19__20_,
         CARRYB_19__19_, CARRYB_19__18_, CARRYB_19__17_, CARRYB_19__16_,
         CARRYB_19__15_, CARRYB_19__14_, CARRYB_19__13_, CARRYB_19__12_,
         CARRYB_19__11_, CARRYB_19__10_, CARRYB_19__9_, CARRYB_19__8_,
         CARRYB_19__7_, CARRYB_19__6_, CARRYB_19__5_, CARRYB_19__4_,
         CARRYB_19__3_, CARRYB_19__2_, CARRYB_19__1_, CARRYB_19__0_,
         CARRYB_18__22_, CARRYB_18__21_, CARRYB_18__20_, CARRYB_18__19_,
         CARRYB_18__18_, CARRYB_18__17_, CARRYB_18__16_, CARRYB_18__15_,
         CARRYB_18__14_, CARRYB_18__13_, CARRYB_18__12_, CARRYB_18__11_,
         CARRYB_18__10_, CARRYB_18__9_, CARRYB_18__8_, CARRYB_18__7_,
         CARRYB_18__6_, CARRYB_18__5_, CARRYB_18__4_, CARRYB_18__3_,
         CARRYB_18__2_, CARRYB_18__1_, CARRYB_18__0_, CARRYB_17__22_,
         CARRYB_17__21_, CARRYB_17__20_, CARRYB_17__19_, CARRYB_17__18_,
         CARRYB_17__17_, CARRYB_17__16_, CARRYB_17__15_, CARRYB_17__14_,
         CARRYB_17__13_, CARRYB_17__12_, CARRYB_17__11_, CARRYB_17__10_,
         CARRYB_17__9_, CARRYB_17__8_, CARRYB_17__7_, CARRYB_17__6_,
         CARRYB_17__5_, CARRYB_17__4_, CARRYB_17__3_, CARRYB_17__2_,
         CARRYB_17__1_, CARRYB_17__0_, CARRYB_16__22_, CARRYB_16__21_,
         CARRYB_16__20_, CARRYB_16__19_, CARRYB_16__18_, CARRYB_16__17_,
         CARRYB_16__16_, CARRYB_16__15_, CARRYB_16__14_, CARRYB_16__13_,
         CARRYB_16__12_, CARRYB_16__11_, CARRYB_16__10_, CARRYB_16__9_,
         CARRYB_16__8_, CARRYB_16__7_, CARRYB_16__6_, CARRYB_16__5_,
         CARRYB_16__4_, CARRYB_16__3_, CARRYB_16__2_, CARRYB_16__1_,
         CARRYB_16__0_, CARRYB_15__22_, CARRYB_15__21_, CARRYB_15__20_,
         CARRYB_15__19_, CARRYB_15__18_, CARRYB_15__17_, CARRYB_15__16_,
         CARRYB_15__15_, CARRYB_15__14_, CARRYB_15__13_, CARRYB_15__12_,
         CARRYB_15__11_, CARRYB_15__10_, CARRYB_15__9_, CARRYB_15__8_,
         CARRYB_15__7_, CARRYB_15__6_, CARRYB_15__5_, CARRYB_15__4_,
         CARRYB_15__3_, CARRYB_15__2_, CARRYB_15__1_, CARRYB_15__0_,
         CARRYB_14__22_, CARRYB_14__21_, CARRYB_14__20_, CARRYB_14__19_,
         CARRYB_14__18_, CARRYB_14__17_, CARRYB_14__16_, CARRYB_14__15_,
         CARRYB_14__14_, CARRYB_14__13_, CARRYB_14__12_, CARRYB_14__11_,
         CARRYB_14__10_, CARRYB_14__9_, CARRYB_14__8_, CARRYB_14__7_,
         CARRYB_14__6_, CARRYB_14__5_, CARRYB_14__4_, CARRYB_14__3_,
         CARRYB_14__2_, CARRYB_14__1_, CARRYB_14__0_, CARRYB_13__22_,
         CARRYB_13__21_, CARRYB_13__20_, CARRYB_13__19_, CARRYB_13__18_,
         CARRYB_13__17_, CARRYB_13__16_, CARRYB_13__15_, CARRYB_13__14_,
         CARRYB_13__13_, CARRYB_13__12_, CARRYB_13__11_, CARRYB_13__10_,
         CARRYB_13__9_, CARRYB_13__8_, CARRYB_13__7_, CARRYB_13__6_,
         CARRYB_13__5_, CARRYB_13__4_, CARRYB_13__3_, CARRYB_13__2_,
         CARRYB_13__1_, CARRYB_13__0_, CARRYB_12__22_, CARRYB_12__21_,
         CARRYB_12__20_, CARRYB_12__19_, CARRYB_12__18_, CARRYB_12__17_,
         CARRYB_12__16_, CARRYB_12__15_, CARRYB_12__14_, CARRYB_12__13_,
         CARRYB_12__12_, CARRYB_12__11_, CARRYB_12__10_, CARRYB_12__9_,
         CARRYB_12__8_, CARRYB_12__7_, CARRYB_12__6_, CARRYB_12__5_,
         CARRYB_12__4_, CARRYB_12__3_, CARRYB_12__2_, CARRYB_12__1_,
         CARRYB_12__0_, CARRYB_11__22_, CARRYB_11__21_, CARRYB_11__20_,
         CARRYB_11__19_, CARRYB_11__18_, CARRYB_11__17_, CARRYB_11__16_,
         CARRYB_11__15_, CARRYB_11__14_, CARRYB_11__13_, CARRYB_11__12_,
         CARRYB_11__11_, CARRYB_11__10_, CARRYB_11__9_, CARRYB_11__8_,
         CARRYB_11__7_, CARRYB_11__6_, CARRYB_11__5_, CARRYB_11__4_,
         CARRYB_11__3_, CARRYB_11__2_, CARRYB_11__1_, CARRYB_11__0_,
         CARRYB_10__22_, CARRYB_10__21_, CARRYB_10__20_, CARRYB_10__19_,
         CARRYB_10__18_, CARRYB_10__17_, CARRYB_10__16_, CARRYB_10__15_,
         CARRYB_10__14_, CARRYB_10__13_, CARRYB_10__12_, CARRYB_10__11_,
         CARRYB_10__10_, CARRYB_10__9_, CARRYB_10__8_, CARRYB_10__7_,
         CARRYB_10__6_, CARRYB_10__5_, CARRYB_10__4_, CARRYB_10__3_,
         CARRYB_10__2_, CARRYB_10__1_, CARRYB_10__0_, CARRYB_9__22_,
         CARRYB_9__21_, CARRYB_9__20_, CARRYB_9__19_, CARRYB_9__18_,
         CARRYB_9__17_, CARRYB_9__16_, CARRYB_9__15_, CARRYB_9__14_,
         CARRYB_9__13_, CARRYB_9__12_, CARRYB_9__11_, CARRYB_9__10_,
         CARRYB_9__9_, CARRYB_9__8_, CARRYB_9__7_, CARRYB_9__6_, CARRYB_9__5_,
         CARRYB_9__4_, CARRYB_9__3_, CARRYB_9__2_, CARRYB_9__1_, CARRYB_9__0_,
         CARRYB_8__22_, CARRYB_8__21_, CARRYB_8__20_, CARRYB_8__19_,
         CARRYB_8__18_, CARRYB_8__17_, CARRYB_8__16_, CARRYB_8__15_,
         CARRYB_8__14_, CARRYB_8__13_, CARRYB_8__12_, CARRYB_8__11_,
         CARRYB_8__10_, CARRYB_8__9_, CARRYB_8__8_, CARRYB_8__7_, CARRYB_8__6_,
         CARRYB_8__5_, CARRYB_8__4_, CARRYB_8__3_, CARRYB_8__2_, CARRYB_8__1_,
         CARRYB_8__0_, CARRYB_7__22_, CARRYB_7__21_, CARRYB_7__20_,
         CARRYB_7__19_, CARRYB_7__18_, CARRYB_7__17_, CARRYB_7__16_,
         CARRYB_7__15_, CARRYB_7__14_, CARRYB_7__13_, CARRYB_7__12_,
         CARRYB_7__11_, CARRYB_7__10_, CARRYB_7__9_, CARRYB_7__8_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__22_,
         CARRYB_6__21_, CARRYB_6__20_, CARRYB_6__19_, CARRYB_6__18_,
         CARRYB_6__17_, CARRYB_6__16_, CARRYB_6__15_, CARRYB_6__14_,
         CARRYB_6__13_, CARRYB_6__12_, CARRYB_6__11_, CARRYB_6__10_,
         CARRYB_6__9_, CARRYB_6__8_, CARRYB_6__7_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__22_, CARRYB_5__21_, CARRYB_5__20_, CARRYB_5__19_,
         CARRYB_5__18_, CARRYB_5__17_, CARRYB_5__16_, CARRYB_5__15_,
         CARRYB_5__14_, CARRYB_5__13_, CARRYB_5__12_, CARRYB_5__11_,
         CARRYB_5__10_, CARRYB_5__9_, CARRYB_5__8_, CARRYB_5__7_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__22_, CARRYB_4__21_, CARRYB_4__20_,
         CARRYB_4__19_, CARRYB_4__18_, CARRYB_4__17_, CARRYB_4__16_,
         CARRYB_4__15_, CARRYB_4__14_, CARRYB_4__13_, CARRYB_4__12_,
         CARRYB_4__11_, CARRYB_4__10_, CARRYB_4__9_, CARRYB_4__8_,
         CARRYB_4__7_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__22_,
         CARRYB_3__21_, CARRYB_3__20_, CARRYB_3__19_, CARRYB_3__18_,
         CARRYB_3__17_, CARRYB_3__16_, CARRYB_3__15_, CARRYB_3__14_,
         CARRYB_3__13_, CARRYB_3__12_, CARRYB_3__11_, CARRYB_3__10_,
         CARRYB_3__9_, CARRYB_3__8_, CARRYB_3__7_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__22_, CARRYB_2__21_, CARRYB_2__20_, CARRYB_2__19_,
         CARRYB_2__18_, CARRYB_2__17_, CARRYB_2__16_, CARRYB_2__15_,
         CARRYB_2__14_, CARRYB_2__13_, CARRYB_2__12_, CARRYB_2__11_,
         CARRYB_2__10_, CARRYB_2__9_, CARRYB_2__8_, CARRYB_2__7_, CARRYB_2__6_,
         CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_, CARRYB_2__1_,
         CARRYB_2__0_, CARRYB_1__0_, SUMB_23__22_, SUMB_23__21_, SUMB_23__20_,
         SUMB_23__19_, SUMB_23__18_, SUMB_23__17_, SUMB_23__16_, SUMB_23__15_,
         SUMB_23__14_, SUMB_23__13_, SUMB_23__12_, SUMB_23__11_, SUMB_23__10_,
         SUMB_23__9_, SUMB_23__8_, SUMB_23__7_, SUMB_23__6_, SUMB_23__5_,
         SUMB_23__4_, SUMB_23__3_, SUMB_23__2_, SUMB_23__1_, SUMB_23__0_,
         SUMB_22__22_, SUMB_22__21_, SUMB_22__20_, SUMB_22__19_, SUMB_22__18_,
         SUMB_22__17_, SUMB_22__16_, SUMB_22__15_, SUMB_22__14_, SUMB_22__13_,
         SUMB_22__12_, SUMB_22__11_, SUMB_22__10_, SUMB_22__9_, SUMB_22__8_,
         SUMB_22__7_, SUMB_22__6_, SUMB_22__5_, SUMB_22__4_, SUMB_22__3_,
         SUMB_22__2_, SUMB_22__1_, SUMB_21__22_, SUMB_21__21_, SUMB_21__20_,
         SUMB_21__19_, SUMB_21__18_, SUMB_21__17_, SUMB_21__16_, SUMB_21__15_,
         SUMB_21__14_, SUMB_21__13_, SUMB_21__12_, SUMB_21__11_, SUMB_21__10_,
         SUMB_21__9_, SUMB_21__8_, SUMB_21__7_, SUMB_21__6_, SUMB_21__5_,
         SUMB_21__4_, SUMB_21__3_, SUMB_21__2_, SUMB_21__1_, SUMB_20__22_,
         SUMB_20__21_, SUMB_20__20_, SUMB_20__19_, SUMB_20__18_, SUMB_20__17_,
         SUMB_20__16_, SUMB_20__15_, SUMB_20__14_, SUMB_20__13_, SUMB_20__12_,
         SUMB_20__11_, SUMB_20__10_, SUMB_20__9_, SUMB_20__8_, SUMB_20__7_,
         SUMB_20__6_, SUMB_20__5_, SUMB_20__4_, SUMB_20__3_, SUMB_20__2_,
         SUMB_20__1_, SUMB_19__22_, SUMB_19__21_, SUMB_19__20_, SUMB_19__19_,
         SUMB_19__18_, SUMB_19__17_, SUMB_19__16_, SUMB_19__15_, SUMB_19__14_,
         SUMB_19__13_, SUMB_19__12_, SUMB_19__11_, SUMB_19__10_, SUMB_19__9_,
         SUMB_19__8_, SUMB_19__7_, SUMB_19__6_, SUMB_19__5_, SUMB_19__4_,
         SUMB_19__3_, SUMB_19__2_, SUMB_19__1_, SUMB_18__22_, SUMB_18__21_,
         SUMB_18__20_, SUMB_18__19_, SUMB_18__18_, SUMB_18__17_, SUMB_18__16_,
         SUMB_18__15_, SUMB_18__14_, SUMB_18__13_, SUMB_18__12_, SUMB_18__11_,
         SUMB_18__10_, SUMB_18__9_, SUMB_18__8_, SUMB_18__7_, SUMB_18__6_,
         SUMB_18__5_, SUMB_18__4_, SUMB_18__3_, SUMB_18__2_, SUMB_18__1_,
         SUMB_17__22_, SUMB_17__21_, SUMB_17__20_, SUMB_17__19_, SUMB_17__18_,
         SUMB_17__17_, SUMB_17__16_, SUMB_17__15_, SUMB_17__14_, SUMB_17__13_,
         SUMB_17__12_, SUMB_17__11_, SUMB_17__10_, SUMB_17__9_, SUMB_17__8_,
         SUMB_17__7_, SUMB_17__6_, SUMB_17__5_, SUMB_17__4_, SUMB_17__3_,
         SUMB_17__2_, SUMB_17__1_, SUMB_16__22_, SUMB_16__21_, SUMB_16__20_,
         SUMB_16__19_, SUMB_16__18_, SUMB_16__17_, SUMB_16__16_, SUMB_16__15_,
         SUMB_16__14_, SUMB_16__13_, SUMB_16__12_, SUMB_16__11_, SUMB_16__10_,
         SUMB_16__9_, SUMB_16__8_, SUMB_16__7_, SUMB_16__6_, SUMB_16__5_,
         SUMB_16__4_, SUMB_16__3_, SUMB_16__2_, SUMB_16__1_, SUMB_15__22_,
         SUMB_15__21_, SUMB_15__20_, SUMB_15__19_, SUMB_15__18_, SUMB_15__17_,
         SUMB_15__16_, SUMB_15__15_, SUMB_15__14_, SUMB_15__13_, SUMB_15__12_,
         SUMB_15__11_, SUMB_15__10_, SUMB_15__9_, SUMB_15__8_, SUMB_15__7_,
         SUMB_15__6_, SUMB_15__5_, SUMB_15__4_, SUMB_15__3_, SUMB_15__2_,
         SUMB_15__1_, SUMB_14__22_, SUMB_14__21_, SUMB_14__20_, SUMB_14__19_,
         SUMB_14__18_, SUMB_14__17_, SUMB_14__16_, SUMB_14__15_, SUMB_14__14_,
         SUMB_14__13_, SUMB_14__12_, SUMB_14__11_, SUMB_14__10_, SUMB_14__9_,
         SUMB_14__8_, SUMB_14__7_, SUMB_14__6_, SUMB_14__5_, SUMB_14__4_,
         SUMB_14__3_, SUMB_14__2_, SUMB_14__1_, SUMB_13__22_, SUMB_13__21_,
         SUMB_13__20_, SUMB_13__19_, SUMB_13__18_, SUMB_13__17_, SUMB_13__16_,
         SUMB_13__15_, SUMB_13__14_, SUMB_13__13_, SUMB_13__12_, SUMB_13__11_,
         SUMB_13__10_, SUMB_13__9_, SUMB_13__8_, SUMB_13__7_, SUMB_13__6_,
         SUMB_13__5_, SUMB_13__4_, SUMB_13__3_, SUMB_13__2_, SUMB_13__1_,
         SUMB_12__22_, SUMB_12__21_, SUMB_12__20_, SUMB_12__19_, SUMB_12__18_,
         SUMB_12__17_, SUMB_12__16_, SUMB_12__15_, SUMB_12__14_, SUMB_12__13_,
         SUMB_12__12_, SUMB_12__11_, SUMB_12__10_, SUMB_12__9_, SUMB_12__8_,
         SUMB_12__7_, SUMB_12__6_, SUMB_12__5_, SUMB_12__4_, SUMB_12__3_,
         SUMB_12__2_, SUMB_12__1_, SUMB_11__22_, SUMB_11__21_, SUMB_11__20_,
         SUMB_11__19_, SUMB_11__18_, SUMB_11__17_, SUMB_11__16_, SUMB_11__15_,
         SUMB_11__14_, SUMB_11__13_, SUMB_11__12_, SUMB_11__11_, SUMB_11__10_,
         SUMB_11__9_, SUMB_11__8_, SUMB_11__7_, SUMB_11__6_, SUMB_11__5_,
         SUMB_11__4_, SUMB_11__3_, SUMB_11__2_, SUMB_11__1_, SUMB_10__22_,
         SUMB_10__21_, SUMB_10__20_, SUMB_10__19_, SUMB_10__18_, SUMB_10__17_,
         SUMB_10__16_, SUMB_10__15_, SUMB_10__14_, SUMB_10__13_, SUMB_10__12_,
         SUMB_10__11_, SUMB_10__10_, SUMB_10__9_, SUMB_10__8_, SUMB_10__7_,
         SUMB_10__6_, SUMB_10__5_, SUMB_10__4_, SUMB_10__3_, SUMB_10__2_,
         SUMB_10__1_, SUMB_9__22_, SUMB_9__21_, SUMB_9__20_, SUMB_9__19_,
         SUMB_9__18_, SUMB_9__17_, SUMB_9__16_, SUMB_9__15_, SUMB_9__14_,
         SUMB_9__13_, SUMB_9__12_, SUMB_9__11_, SUMB_9__10_, SUMB_9__9_,
         SUMB_9__8_, SUMB_9__7_, SUMB_9__6_, SUMB_9__5_, SUMB_9__4_,
         SUMB_9__3_, SUMB_9__2_, SUMB_9__1_, SUMB_8__22_, SUMB_8__21_,
         SUMB_8__20_, SUMB_8__19_, SUMB_8__18_, SUMB_8__17_, SUMB_8__16_,
         SUMB_8__15_, SUMB_8__14_, SUMB_8__13_, SUMB_8__12_, SUMB_8__11_,
         SUMB_8__10_, SUMB_8__9_, SUMB_8__8_, SUMB_8__7_, SUMB_8__6_,
         SUMB_8__5_, SUMB_8__4_, SUMB_8__3_, SUMB_8__2_, SUMB_8__1_,
         SUMB_7__22_, SUMB_7__21_, SUMB_7__20_, SUMB_7__19_, SUMB_7__18_,
         SUMB_7__17_, SUMB_7__16_, SUMB_7__15_, SUMB_7__14_, SUMB_7__13_,
         SUMB_7__12_, SUMB_7__11_, SUMB_7__10_, SUMB_7__9_, SUMB_7__8_,
         SUMB_7__7_, SUMB_7__6_, SUMB_7__5_, SUMB_7__4_, SUMB_7__3_,
         SUMB_7__2_, SUMB_7__1_, SUMB_6__22_, SUMB_6__21_, SUMB_6__20_,
         SUMB_6__19_, SUMB_6__18_, SUMB_6__17_, SUMB_6__16_, SUMB_6__15_,
         SUMB_6__14_, SUMB_6__13_, SUMB_6__12_, SUMB_6__11_, SUMB_6__10_,
         SUMB_6__9_, SUMB_6__8_, SUMB_6__7_, SUMB_6__6_, SUMB_6__5_,
         SUMB_6__4_, SUMB_6__3_, SUMB_6__2_, SUMB_6__1_, SUMB_5__22_,
         SUMB_5__21_, SUMB_5__20_, SUMB_5__19_, SUMB_5__18_, SUMB_5__17_,
         SUMB_5__16_, SUMB_5__15_, SUMB_5__14_, SUMB_5__13_, SUMB_5__12_,
         SUMB_5__11_, SUMB_5__10_, SUMB_5__9_, SUMB_5__8_, SUMB_5__7_,
         SUMB_5__6_, SUMB_5__5_, SUMB_5__4_, SUMB_5__3_, SUMB_5__2_,
         SUMB_5__1_, SUMB_4__22_, SUMB_4__21_, SUMB_4__20_, SUMB_4__19_,
         SUMB_4__18_, SUMB_4__17_, SUMB_4__16_, SUMB_4__15_, SUMB_4__14_,
         SUMB_4__13_, SUMB_4__12_, SUMB_4__11_, SUMB_4__10_, SUMB_4__9_,
         SUMB_4__8_, SUMB_4__7_, SUMB_4__6_, SUMB_4__5_, SUMB_4__4_,
         SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__22_, SUMB_3__21_,
         SUMB_3__20_, SUMB_3__19_, SUMB_3__18_, SUMB_3__17_, SUMB_3__16_,
         SUMB_3__15_, SUMB_3__14_, SUMB_3__13_, SUMB_3__12_, SUMB_3__11_,
         SUMB_3__10_, SUMB_3__9_, SUMB_3__8_, SUMB_3__7_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__22_, SUMB_2__21_, SUMB_2__20_, SUMB_2__19_, SUMB_2__18_,
         SUMB_2__17_, SUMB_2__16_, SUMB_2__15_, SUMB_2__14_, SUMB_2__13_,
         SUMB_2__12_, SUMB_2__11_, SUMB_2__10_, SUMB_2__9_, SUMB_2__8_,
         SUMB_2__7_, SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_,
         SUMB_2__2_, SUMB_2__1_, A1_20_, A1_19_, A1_18_, A1_17_, A1_16_,
         A1_15_, A1_14_, A1_13_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21;

  FA_X1 S4_0 ( .A(ab_23__0_), .B(CARRYB_22__0_), .CI(SUMB_22__1_), .CO(
        CARRYB_23__0_), .S(SUMB_23__0_) );
  FA_X1 S4_1 ( .A(ab_23__1_), .B(CARRYB_22__1_), .CI(SUMB_22__2_), .CO(
        CARRYB_23__1_), .S(SUMB_23__1_) );
  FA_X1 S4_2 ( .A(ab_23__2_), .B(CARRYB_22__2_), .CI(SUMB_22__3_), .CO(
        CARRYB_23__2_), .S(SUMB_23__2_) );
  FA_X1 S4_3 ( .A(ab_23__3_), .B(CARRYB_22__3_), .CI(SUMB_22__4_), .CO(
        CARRYB_23__3_), .S(SUMB_23__3_) );
  FA_X1 S4_4 ( .A(ab_23__4_), .B(CARRYB_22__4_), .CI(SUMB_22__5_), .CO(
        CARRYB_23__4_), .S(SUMB_23__4_) );
  FA_X1 S4_5 ( .A(ab_23__5_), .B(CARRYB_22__5_), .CI(SUMB_22__6_), .CO(
        CARRYB_23__5_), .S(SUMB_23__5_) );
  FA_X1 S4_6 ( .A(ab_23__6_), .B(CARRYB_22__6_), .CI(SUMB_22__7_), .CO(
        CARRYB_23__6_), .S(SUMB_23__6_) );
  FA_X1 S4_7 ( .A(ab_23__7_), .B(CARRYB_22__7_), .CI(SUMB_22__8_), .CO(
        CARRYB_23__7_), .S(SUMB_23__7_) );
  FA_X1 S4_8 ( .A(ab_23__8_), .B(CARRYB_22__8_), .CI(SUMB_22__9_), .CO(
        CARRYB_23__8_), .S(SUMB_23__8_) );
  FA_X1 S4_9 ( .A(ab_23__9_), .B(CARRYB_22__9_), .CI(SUMB_22__10_), .CO(
        CARRYB_23__9_), .S(SUMB_23__9_) );
  FA_X1 S4_10 ( .A(ab_23__10_), .B(CARRYB_22__10_), .CI(SUMB_22__11_), .CO(
        CARRYB_23__10_), .S(SUMB_23__10_) );
  FA_X1 S4_11 ( .A(ab_23__11_), .B(CARRYB_22__11_), .CI(SUMB_22__12_), .CO(
        CARRYB_23__11_), .S(SUMB_23__11_) );
  FA_X1 S4_12 ( .A(ab_23__12_), .B(CARRYB_22__12_), .CI(SUMB_22__13_), .CO(
        CARRYB_23__12_), .S(SUMB_23__12_) );
  FA_X1 S4_13 ( .A(ab_23__13_), .B(CARRYB_22__13_), .CI(SUMB_22__14_), .CO(
        CARRYB_23__13_), .S(SUMB_23__13_) );
  FA_X1 S4_14 ( .A(ab_23__14_), .B(CARRYB_22__14_), .CI(SUMB_22__15_), .CO(
        CARRYB_23__14_), .S(SUMB_23__14_) );
  FA_X1 S4_15 ( .A(ab_23__15_), .B(CARRYB_22__15_), .CI(SUMB_22__16_), .CO(
        CARRYB_23__15_), .S(SUMB_23__15_) );
  FA_X1 S4_16 ( .A(ab_23__16_), .B(CARRYB_22__16_), .CI(SUMB_22__17_), .CO(
        CARRYB_23__16_), .S(SUMB_23__16_) );
  FA_X1 S4_17 ( .A(ab_23__17_), .B(CARRYB_22__17_), .CI(SUMB_22__18_), .CO(
        CARRYB_23__17_), .S(SUMB_23__17_) );
  FA_X1 S4_18 ( .A(ab_23__18_), .B(CARRYB_22__18_), .CI(SUMB_22__19_), .CO(
        CARRYB_23__18_), .S(SUMB_23__18_) );
  FA_X1 S4_19 ( .A(ab_23__19_), .B(CARRYB_22__19_), .CI(SUMB_22__20_), .CO(
        CARRYB_23__19_), .S(SUMB_23__19_) );
  FA_X1 S4_20 ( .A(ab_23__20_), .B(CARRYB_22__20_), .CI(SUMB_22__21_), .CO(
        CARRYB_23__20_), .S(SUMB_23__20_) );
  FA_X1 S4_21 ( .A(ab_23__21_), .B(CARRYB_22__21_), .CI(SUMB_22__22_), .CO(
        CARRYB_23__21_), .S(SUMB_23__21_) );
  FA_X1 S5_22 ( .A(ab_23__22_), .B(CARRYB_22__22_), .CI(ab_22__23_), .CO(
        CARRYB_23__22_), .S(SUMB_23__22_) );
  FA_X1 S1_22_0 ( .A(ab_22__0_), .B(CARRYB_21__0_), .CI(SUMB_21__1_), .CO(
        CARRYB_22__0_), .S(A1_20_) );
  FA_X1 S2_22_1 ( .A(ab_22__1_), .B(CARRYB_21__1_), .CI(SUMB_21__2_), .CO(
        CARRYB_22__1_), .S(SUMB_22__1_) );
  FA_X1 S2_22_2 ( .A(ab_22__2_), .B(CARRYB_21__2_), .CI(SUMB_21__3_), .CO(
        CARRYB_22__2_), .S(SUMB_22__2_) );
  FA_X1 S2_22_3 ( .A(ab_22__3_), .B(CARRYB_21__3_), .CI(SUMB_21__4_), .CO(
        CARRYB_22__3_), .S(SUMB_22__3_) );
  FA_X1 S2_22_4 ( .A(ab_22__4_), .B(CARRYB_21__4_), .CI(SUMB_21__5_), .CO(
        CARRYB_22__4_), .S(SUMB_22__4_) );
  FA_X1 S2_22_5 ( .A(ab_22__5_), .B(CARRYB_21__5_), .CI(SUMB_21__6_), .CO(
        CARRYB_22__5_), .S(SUMB_22__5_) );
  FA_X1 S2_22_6 ( .A(ab_22__6_), .B(CARRYB_21__6_), .CI(SUMB_21__7_), .CO(
        CARRYB_22__6_), .S(SUMB_22__6_) );
  FA_X1 S2_22_7 ( .A(ab_22__7_), .B(CARRYB_21__7_), .CI(SUMB_21__8_), .CO(
        CARRYB_22__7_), .S(SUMB_22__7_) );
  FA_X1 S2_22_8 ( .A(ab_22__8_), .B(CARRYB_21__8_), .CI(SUMB_21__9_), .CO(
        CARRYB_22__8_), .S(SUMB_22__8_) );
  FA_X1 S2_22_9 ( .A(ab_22__9_), .B(CARRYB_21__9_), .CI(SUMB_21__10_), .CO(
        CARRYB_22__9_), .S(SUMB_22__9_) );
  FA_X1 S2_22_10 ( .A(ab_22__10_), .B(CARRYB_21__10_), .CI(SUMB_21__11_), .CO(
        CARRYB_22__10_), .S(SUMB_22__10_) );
  FA_X1 S2_22_11 ( .A(ab_22__11_), .B(CARRYB_21__11_), .CI(SUMB_21__12_), .CO(
        CARRYB_22__11_), .S(SUMB_22__11_) );
  FA_X1 S2_22_12 ( .A(ab_22__12_), .B(CARRYB_21__12_), .CI(SUMB_21__13_), .CO(
        CARRYB_22__12_), .S(SUMB_22__12_) );
  FA_X1 S2_22_13 ( .A(ab_22__13_), .B(CARRYB_21__13_), .CI(SUMB_21__14_), .CO(
        CARRYB_22__13_), .S(SUMB_22__13_) );
  FA_X1 S2_22_14 ( .A(ab_22__14_), .B(CARRYB_21__14_), .CI(SUMB_21__15_), .CO(
        CARRYB_22__14_), .S(SUMB_22__14_) );
  FA_X1 S2_22_15 ( .A(ab_22__15_), .B(CARRYB_21__15_), .CI(SUMB_21__16_), .CO(
        CARRYB_22__15_), .S(SUMB_22__15_) );
  FA_X1 S2_22_16 ( .A(ab_22__16_), .B(CARRYB_21__16_), .CI(SUMB_21__17_), .CO(
        CARRYB_22__16_), .S(SUMB_22__16_) );
  FA_X1 S2_22_17 ( .A(ab_22__17_), .B(CARRYB_21__17_), .CI(SUMB_21__18_), .CO(
        CARRYB_22__17_), .S(SUMB_22__17_) );
  FA_X1 S2_22_18 ( .A(ab_22__18_), .B(CARRYB_21__18_), .CI(SUMB_21__19_), .CO(
        CARRYB_22__18_), .S(SUMB_22__18_) );
  FA_X1 S2_22_19 ( .A(ab_22__19_), .B(CARRYB_21__19_), .CI(SUMB_21__20_), .CO(
        CARRYB_22__19_), .S(SUMB_22__19_) );
  FA_X1 S2_22_20 ( .A(ab_22__20_), .B(CARRYB_21__20_), .CI(SUMB_21__21_), .CO(
        CARRYB_22__20_), .S(SUMB_22__20_) );
  FA_X1 S2_22_21 ( .A(ab_22__21_), .B(CARRYB_21__21_), .CI(SUMB_21__22_), .CO(
        CARRYB_22__21_), .S(SUMB_22__21_) );
  FA_X1 S3_22_22 ( .A(ab_22__22_), .B(CARRYB_21__22_), .CI(ab_21__23_), .CO(
        CARRYB_22__22_), .S(SUMB_22__22_) );
  FA_X1 S1_21_0 ( .A(ab_21__0_), .B(CARRYB_20__0_), .CI(SUMB_20__1_), .CO(
        CARRYB_21__0_), .S(A1_19_) );
  FA_X1 S2_21_1 ( .A(ab_21__1_), .B(CARRYB_20__1_), .CI(SUMB_20__2_), .CO(
        CARRYB_21__1_), .S(SUMB_21__1_) );
  FA_X1 S2_21_2 ( .A(ab_21__2_), .B(CARRYB_20__2_), .CI(SUMB_20__3_), .CO(
        CARRYB_21__2_), .S(SUMB_21__2_) );
  FA_X1 S2_21_3 ( .A(ab_21__3_), .B(CARRYB_20__3_), .CI(SUMB_20__4_), .CO(
        CARRYB_21__3_), .S(SUMB_21__3_) );
  FA_X1 S2_21_4 ( .A(ab_21__4_), .B(CARRYB_20__4_), .CI(SUMB_20__5_), .CO(
        CARRYB_21__4_), .S(SUMB_21__4_) );
  FA_X1 S2_21_5 ( .A(ab_21__5_), .B(CARRYB_20__5_), .CI(SUMB_20__6_), .CO(
        CARRYB_21__5_), .S(SUMB_21__5_) );
  FA_X1 S2_21_6 ( .A(ab_21__6_), .B(CARRYB_20__6_), .CI(SUMB_20__7_), .CO(
        CARRYB_21__6_), .S(SUMB_21__6_) );
  FA_X1 S2_21_7 ( .A(ab_21__7_), .B(CARRYB_20__7_), .CI(SUMB_20__8_), .CO(
        CARRYB_21__7_), .S(SUMB_21__7_) );
  FA_X1 S2_21_8 ( .A(ab_21__8_), .B(CARRYB_20__8_), .CI(SUMB_20__9_), .CO(
        CARRYB_21__8_), .S(SUMB_21__8_) );
  FA_X1 S2_21_9 ( .A(ab_21__9_), .B(CARRYB_20__9_), .CI(SUMB_20__10_), .CO(
        CARRYB_21__9_), .S(SUMB_21__9_) );
  FA_X1 S2_21_10 ( .A(ab_21__10_), .B(CARRYB_20__10_), .CI(SUMB_20__11_), .CO(
        CARRYB_21__10_), .S(SUMB_21__10_) );
  FA_X1 S2_21_11 ( .A(ab_21__11_), .B(CARRYB_20__11_), .CI(SUMB_20__12_), .CO(
        CARRYB_21__11_), .S(SUMB_21__11_) );
  FA_X1 S2_21_12 ( .A(ab_21__12_), .B(CARRYB_20__12_), .CI(SUMB_20__13_), .CO(
        CARRYB_21__12_), .S(SUMB_21__12_) );
  FA_X1 S2_21_13 ( .A(ab_21__13_), .B(CARRYB_20__13_), .CI(SUMB_20__14_), .CO(
        CARRYB_21__13_), .S(SUMB_21__13_) );
  FA_X1 S2_21_14 ( .A(ab_21__14_), .B(CARRYB_20__14_), .CI(SUMB_20__15_), .CO(
        CARRYB_21__14_), .S(SUMB_21__14_) );
  FA_X1 S2_21_15 ( .A(ab_21__15_), .B(CARRYB_20__15_), .CI(SUMB_20__16_), .CO(
        CARRYB_21__15_), .S(SUMB_21__15_) );
  FA_X1 S2_21_16 ( .A(ab_21__16_), .B(CARRYB_20__16_), .CI(SUMB_20__17_), .CO(
        CARRYB_21__16_), .S(SUMB_21__16_) );
  FA_X1 S2_21_17 ( .A(ab_21__17_), .B(CARRYB_20__17_), .CI(SUMB_20__18_), .CO(
        CARRYB_21__17_), .S(SUMB_21__17_) );
  FA_X1 S2_21_18 ( .A(ab_21__18_), .B(CARRYB_20__18_), .CI(SUMB_20__19_), .CO(
        CARRYB_21__18_), .S(SUMB_21__18_) );
  FA_X1 S2_21_19 ( .A(ab_21__19_), .B(CARRYB_20__19_), .CI(SUMB_20__20_), .CO(
        CARRYB_21__19_), .S(SUMB_21__19_) );
  FA_X1 S2_21_20 ( .A(ab_21__20_), .B(CARRYB_20__20_), .CI(SUMB_20__21_), .CO(
        CARRYB_21__20_), .S(SUMB_21__20_) );
  FA_X1 S2_21_21 ( .A(ab_21__21_), .B(CARRYB_20__21_), .CI(SUMB_20__22_), .CO(
        CARRYB_21__21_), .S(SUMB_21__21_) );
  FA_X1 S3_21_22 ( .A(ab_21__22_), .B(CARRYB_20__22_), .CI(ab_20__23_), .CO(
        CARRYB_21__22_), .S(SUMB_21__22_) );
  FA_X1 S1_20_0 ( .A(ab_20__0_), .B(CARRYB_19__0_), .CI(SUMB_19__1_), .CO(
        CARRYB_20__0_), .S(A1_18_) );
  FA_X1 S2_20_1 ( .A(ab_20__1_), .B(CARRYB_19__1_), .CI(SUMB_19__2_), .CO(
        CARRYB_20__1_), .S(SUMB_20__1_) );
  FA_X1 S2_20_2 ( .A(ab_20__2_), .B(CARRYB_19__2_), .CI(SUMB_19__3_), .CO(
        CARRYB_20__2_), .S(SUMB_20__2_) );
  FA_X1 S2_20_3 ( .A(ab_20__3_), .B(CARRYB_19__3_), .CI(SUMB_19__4_), .CO(
        CARRYB_20__3_), .S(SUMB_20__3_) );
  FA_X1 S2_20_4 ( .A(ab_20__4_), .B(CARRYB_19__4_), .CI(SUMB_19__5_), .CO(
        CARRYB_20__4_), .S(SUMB_20__4_) );
  FA_X1 S2_20_5 ( .A(ab_20__5_), .B(CARRYB_19__5_), .CI(SUMB_19__6_), .CO(
        CARRYB_20__5_), .S(SUMB_20__5_) );
  FA_X1 S2_20_6 ( .A(ab_20__6_), .B(CARRYB_19__6_), .CI(SUMB_19__7_), .CO(
        CARRYB_20__6_), .S(SUMB_20__6_) );
  FA_X1 S2_20_7 ( .A(ab_20__7_), .B(CARRYB_19__7_), .CI(SUMB_19__8_), .CO(
        CARRYB_20__7_), .S(SUMB_20__7_) );
  FA_X1 S2_20_8 ( .A(ab_20__8_), .B(CARRYB_19__8_), .CI(SUMB_19__9_), .CO(
        CARRYB_20__8_), .S(SUMB_20__8_) );
  FA_X1 S2_20_9 ( .A(ab_20__9_), .B(CARRYB_19__9_), .CI(SUMB_19__10_), .CO(
        CARRYB_20__9_), .S(SUMB_20__9_) );
  FA_X1 S2_20_10 ( .A(ab_20__10_), .B(CARRYB_19__10_), .CI(SUMB_19__11_), .CO(
        CARRYB_20__10_), .S(SUMB_20__10_) );
  FA_X1 S2_20_11 ( .A(ab_20__11_), .B(CARRYB_19__11_), .CI(SUMB_19__12_), .CO(
        CARRYB_20__11_), .S(SUMB_20__11_) );
  FA_X1 S2_20_12 ( .A(ab_20__12_), .B(CARRYB_19__12_), .CI(SUMB_19__13_), .CO(
        CARRYB_20__12_), .S(SUMB_20__12_) );
  FA_X1 S2_20_13 ( .A(ab_20__13_), .B(CARRYB_19__13_), .CI(SUMB_19__14_), .CO(
        CARRYB_20__13_), .S(SUMB_20__13_) );
  FA_X1 S2_20_14 ( .A(ab_20__14_), .B(CARRYB_19__14_), .CI(SUMB_19__15_), .CO(
        CARRYB_20__14_), .S(SUMB_20__14_) );
  FA_X1 S2_20_15 ( .A(ab_20__15_), .B(CARRYB_19__15_), .CI(SUMB_19__16_), .CO(
        CARRYB_20__15_), .S(SUMB_20__15_) );
  FA_X1 S2_20_16 ( .A(ab_20__16_), .B(CARRYB_19__16_), .CI(SUMB_19__17_), .CO(
        CARRYB_20__16_), .S(SUMB_20__16_) );
  FA_X1 S2_20_17 ( .A(ab_20__17_), .B(CARRYB_19__17_), .CI(SUMB_19__18_), .CO(
        CARRYB_20__17_), .S(SUMB_20__17_) );
  FA_X1 S2_20_18 ( .A(ab_20__18_), .B(CARRYB_19__18_), .CI(SUMB_19__19_), .CO(
        CARRYB_20__18_), .S(SUMB_20__18_) );
  FA_X1 S2_20_19 ( .A(ab_20__19_), .B(CARRYB_19__19_), .CI(SUMB_19__20_), .CO(
        CARRYB_20__19_), .S(SUMB_20__19_) );
  FA_X1 S2_20_20 ( .A(ab_20__20_), .B(CARRYB_19__20_), .CI(SUMB_19__21_), .CO(
        CARRYB_20__20_), .S(SUMB_20__20_) );
  FA_X1 S2_20_21 ( .A(ab_20__21_), .B(CARRYB_19__21_), .CI(SUMB_19__22_), .CO(
        CARRYB_20__21_), .S(SUMB_20__21_) );
  FA_X1 S3_20_22 ( .A(ab_20__22_), .B(CARRYB_19__22_), .CI(ab_19__23_), .CO(
        CARRYB_20__22_), .S(SUMB_20__22_) );
  FA_X1 S1_19_0 ( .A(ab_19__0_), .B(CARRYB_18__0_), .CI(SUMB_18__1_), .CO(
        CARRYB_19__0_), .S(A1_17_) );
  FA_X1 S2_19_1 ( .A(ab_19__1_), .B(CARRYB_18__1_), .CI(SUMB_18__2_), .CO(
        CARRYB_19__1_), .S(SUMB_19__1_) );
  FA_X1 S2_19_2 ( .A(ab_19__2_), .B(CARRYB_18__2_), .CI(SUMB_18__3_), .CO(
        CARRYB_19__2_), .S(SUMB_19__2_) );
  FA_X1 S2_19_3 ( .A(ab_19__3_), .B(CARRYB_18__3_), .CI(SUMB_18__4_), .CO(
        CARRYB_19__3_), .S(SUMB_19__3_) );
  FA_X1 S2_19_4 ( .A(ab_19__4_), .B(CARRYB_18__4_), .CI(SUMB_18__5_), .CO(
        CARRYB_19__4_), .S(SUMB_19__4_) );
  FA_X1 S2_19_5 ( .A(ab_19__5_), .B(CARRYB_18__5_), .CI(SUMB_18__6_), .CO(
        CARRYB_19__5_), .S(SUMB_19__5_) );
  FA_X1 S2_19_6 ( .A(ab_19__6_), .B(CARRYB_18__6_), .CI(SUMB_18__7_), .CO(
        CARRYB_19__6_), .S(SUMB_19__6_) );
  FA_X1 S2_19_7 ( .A(ab_19__7_), .B(CARRYB_18__7_), .CI(SUMB_18__8_), .CO(
        CARRYB_19__7_), .S(SUMB_19__7_) );
  FA_X1 S2_19_8 ( .A(ab_19__8_), .B(CARRYB_18__8_), .CI(SUMB_18__9_), .CO(
        CARRYB_19__8_), .S(SUMB_19__8_) );
  FA_X1 S2_19_9 ( .A(ab_19__9_), .B(CARRYB_18__9_), .CI(SUMB_18__10_), .CO(
        CARRYB_19__9_), .S(SUMB_19__9_) );
  FA_X1 S2_19_10 ( .A(ab_19__10_), .B(CARRYB_18__10_), .CI(SUMB_18__11_), .CO(
        CARRYB_19__10_), .S(SUMB_19__10_) );
  FA_X1 S2_19_11 ( .A(ab_19__11_), .B(CARRYB_18__11_), .CI(SUMB_18__12_), .CO(
        CARRYB_19__11_), .S(SUMB_19__11_) );
  FA_X1 S2_19_12 ( .A(ab_19__12_), .B(CARRYB_18__12_), .CI(SUMB_18__13_), .CO(
        CARRYB_19__12_), .S(SUMB_19__12_) );
  FA_X1 S2_19_13 ( .A(ab_19__13_), .B(CARRYB_18__13_), .CI(SUMB_18__14_), .CO(
        CARRYB_19__13_), .S(SUMB_19__13_) );
  FA_X1 S2_19_14 ( .A(ab_19__14_), .B(CARRYB_18__14_), .CI(SUMB_18__15_), .CO(
        CARRYB_19__14_), .S(SUMB_19__14_) );
  FA_X1 S2_19_15 ( .A(ab_19__15_), .B(CARRYB_18__15_), .CI(SUMB_18__16_), .CO(
        CARRYB_19__15_), .S(SUMB_19__15_) );
  FA_X1 S2_19_16 ( .A(ab_19__16_), .B(CARRYB_18__16_), .CI(SUMB_18__17_), .CO(
        CARRYB_19__16_), .S(SUMB_19__16_) );
  FA_X1 S2_19_17 ( .A(ab_19__17_), .B(CARRYB_18__17_), .CI(SUMB_18__18_), .CO(
        CARRYB_19__17_), .S(SUMB_19__17_) );
  FA_X1 S2_19_18 ( .A(ab_19__18_), .B(CARRYB_18__18_), .CI(SUMB_18__19_), .CO(
        CARRYB_19__18_), .S(SUMB_19__18_) );
  FA_X1 S2_19_19 ( .A(ab_19__19_), .B(CARRYB_18__19_), .CI(SUMB_18__20_), .CO(
        CARRYB_19__19_), .S(SUMB_19__19_) );
  FA_X1 S2_19_20 ( .A(ab_19__20_), .B(CARRYB_18__20_), .CI(SUMB_18__21_), .CO(
        CARRYB_19__20_), .S(SUMB_19__20_) );
  FA_X1 S2_19_21 ( .A(ab_19__21_), .B(CARRYB_18__21_), .CI(SUMB_18__22_), .CO(
        CARRYB_19__21_), .S(SUMB_19__21_) );
  FA_X1 S3_19_22 ( .A(ab_19__22_), .B(CARRYB_18__22_), .CI(ab_18__23_), .CO(
        CARRYB_19__22_), .S(SUMB_19__22_) );
  FA_X1 S1_18_0 ( .A(ab_18__0_), .B(CARRYB_17__0_), .CI(SUMB_17__1_), .CO(
        CARRYB_18__0_), .S(A1_16_) );
  FA_X1 S2_18_1 ( .A(ab_18__1_), .B(CARRYB_17__1_), .CI(SUMB_17__2_), .CO(
        CARRYB_18__1_), .S(SUMB_18__1_) );
  FA_X1 S2_18_2 ( .A(ab_18__2_), .B(CARRYB_17__2_), .CI(SUMB_17__3_), .CO(
        CARRYB_18__2_), .S(SUMB_18__2_) );
  FA_X1 S2_18_3 ( .A(ab_18__3_), .B(CARRYB_17__3_), .CI(SUMB_17__4_), .CO(
        CARRYB_18__3_), .S(SUMB_18__3_) );
  FA_X1 S2_18_4 ( .A(ab_18__4_), .B(CARRYB_17__4_), .CI(SUMB_17__5_), .CO(
        CARRYB_18__4_), .S(SUMB_18__4_) );
  FA_X1 S2_18_5 ( .A(ab_18__5_), .B(CARRYB_17__5_), .CI(SUMB_17__6_), .CO(
        CARRYB_18__5_), .S(SUMB_18__5_) );
  FA_X1 S2_18_6 ( .A(ab_18__6_), .B(CARRYB_17__6_), .CI(SUMB_17__7_), .CO(
        CARRYB_18__6_), .S(SUMB_18__6_) );
  FA_X1 S2_18_7 ( .A(ab_18__7_), .B(CARRYB_17__7_), .CI(SUMB_17__8_), .CO(
        CARRYB_18__7_), .S(SUMB_18__7_) );
  FA_X1 S2_18_8 ( .A(ab_18__8_), .B(CARRYB_17__8_), .CI(SUMB_17__9_), .CO(
        CARRYB_18__8_), .S(SUMB_18__8_) );
  FA_X1 S2_18_9 ( .A(ab_18__9_), .B(CARRYB_17__9_), .CI(SUMB_17__10_), .CO(
        CARRYB_18__9_), .S(SUMB_18__9_) );
  FA_X1 S2_18_10 ( .A(ab_18__10_), .B(CARRYB_17__10_), .CI(SUMB_17__11_), .CO(
        CARRYB_18__10_), .S(SUMB_18__10_) );
  FA_X1 S2_18_11 ( .A(ab_18__11_), .B(CARRYB_17__11_), .CI(SUMB_17__12_), .CO(
        CARRYB_18__11_), .S(SUMB_18__11_) );
  FA_X1 S2_18_12 ( .A(ab_18__12_), .B(CARRYB_17__12_), .CI(SUMB_17__13_), .CO(
        CARRYB_18__12_), .S(SUMB_18__12_) );
  FA_X1 S2_18_13 ( .A(ab_18__13_), .B(CARRYB_17__13_), .CI(SUMB_17__14_), .CO(
        CARRYB_18__13_), .S(SUMB_18__13_) );
  FA_X1 S2_18_14 ( .A(ab_18__14_), .B(CARRYB_17__14_), .CI(SUMB_17__15_), .CO(
        CARRYB_18__14_), .S(SUMB_18__14_) );
  FA_X1 S2_18_15 ( .A(ab_18__15_), .B(CARRYB_17__15_), .CI(SUMB_17__16_), .CO(
        CARRYB_18__15_), .S(SUMB_18__15_) );
  FA_X1 S2_18_16 ( .A(ab_18__16_), .B(CARRYB_17__16_), .CI(SUMB_17__17_), .CO(
        CARRYB_18__16_), .S(SUMB_18__16_) );
  FA_X1 S2_18_17 ( .A(ab_18__17_), .B(CARRYB_17__17_), .CI(SUMB_17__18_), .CO(
        CARRYB_18__17_), .S(SUMB_18__17_) );
  FA_X1 S2_18_18 ( .A(ab_18__18_), .B(CARRYB_17__18_), .CI(SUMB_17__19_), .CO(
        CARRYB_18__18_), .S(SUMB_18__18_) );
  FA_X1 S2_18_19 ( .A(ab_18__19_), .B(CARRYB_17__19_), .CI(SUMB_17__20_), .CO(
        CARRYB_18__19_), .S(SUMB_18__19_) );
  FA_X1 S2_18_20 ( .A(ab_18__20_), .B(CARRYB_17__20_), .CI(SUMB_17__21_), .CO(
        CARRYB_18__20_), .S(SUMB_18__20_) );
  FA_X1 S2_18_21 ( .A(ab_18__21_), .B(CARRYB_17__21_), .CI(SUMB_17__22_), .CO(
        CARRYB_18__21_), .S(SUMB_18__21_) );
  FA_X1 S3_18_22 ( .A(ab_18__22_), .B(CARRYB_17__22_), .CI(ab_17__23_), .CO(
        CARRYB_18__22_), .S(SUMB_18__22_) );
  FA_X1 S1_17_0 ( .A(ab_17__0_), .B(CARRYB_16__0_), .CI(SUMB_16__1_), .CO(
        CARRYB_17__0_), .S(A1_15_) );
  FA_X1 S2_17_1 ( .A(ab_17__1_), .B(CARRYB_16__1_), .CI(SUMB_16__2_), .CO(
        CARRYB_17__1_), .S(SUMB_17__1_) );
  FA_X1 S2_17_2 ( .A(ab_17__2_), .B(CARRYB_16__2_), .CI(SUMB_16__3_), .CO(
        CARRYB_17__2_), .S(SUMB_17__2_) );
  FA_X1 S2_17_3 ( .A(ab_17__3_), .B(CARRYB_16__3_), .CI(SUMB_16__4_), .CO(
        CARRYB_17__3_), .S(SUMB_17__3_) );
  FA_X1 S2_17_4 ( .A(ab_17__4_), .B(CARRYB_16__4_), .CI(SUMB_16__5_), .CO(
        CARRYB_17__4_), .S(SUMB_17__4_) );
  FA_X1 S2_17_5 ( .A(ab_17__5_), .B(CARRYB_16__5_), .CI(SUMB_16__6_), .CO(
        CARRYB_17__5_), .S(SUMB_17__5_) );
  FA_X1 S2_17_6 ( .A(ab_17__6_), .B(CARRYB_16__6_), .CI(SUMB_16__7_), .CO(
        CARRYB_17__6_), .S(SUMB_17__6_) );
  FA_X1 S2_17_7 ( .A(ab_17__7_), .B(CARRYB_16__7_), .CI(SUMB_16__8_), .CO(
        CARRYB_17__7_), .S(SUMB_17__7_) );
  FA_X1 S2_17_8 ( .A(ab_17__8_), .B(CARRYB_16__8_), .CI(SUMB_16__9_), .CO(
        CARRYB_17__8_), .S(SUMB_17__8_) );
  FA_X1 S2_17_9 ( .A(ab_17__9_), .B(CARRYB_16__9_), .CI(SUMB_16__10_), .CO(
        CARRYB_17__9_), .S(SUMB_17__9_) );
  FA_X1 S2_17_10 ( .A(ab_17__10_), .B(CARRYB_16__10_), .CI(SUMB_16__11_), .CO(
        CARRYB_17__10_), .S(SUMB_17__10_) );
  FA_X1 S2_17_11 ( .A(ab_17__11_), .B(CARRYB_16__11_), .CI(SUMB_16__12_), .CO(
        CARRYB_17__11_), .S(SUMB_17__11_) );
  FA_X1 S2_17_12 ( .A(ab_17__12_), .B(CARRYB_16__12_), .CI(SUMB_16__13_), .CO(
        CARRYB_17__12_), .S(SUMB_17__12_) );
  FA_X1 S2_17_13 ( .A(ab_17__13_), .B(CARRYB_16__13_), .CI(SUMB_16__14_), .CO(
        CARRYB_17__13_), .S(SUMB_17__13_) );
  FA_X1 S2_17_14 ( .A(ab_17__14_), .B(CARRYB_16__14_), .CI(SUMB_16__15_), .CO(
        CARRYB_17__14_), .S(SUMB_17__14_) );
  FA_X1 S2_17_15 ( .A(ab_17__15_), .B(CARRYB_16__15_), .CI(SUMB_16__16_), .CO(
        CARRYB_17__15_), .S(SUMB_17__15_) );
  FA_X1 S2_17_16 ( .A(ab_17__16_), .B(CARRYB_16__16_), .CI(SUMB_16__17_), .CO(
        CARRYB_17__16_), .S(SUMB_17__16_) );
  FA_X1 S2_17_17 ( .A(ab_17__17_), .B(CARRYB_16__17_), .CI(SUMB_16__18_), .CO(
        CARRYB_17__17_), .S(SUMB_17__17_) );
  FA_X1 S2_17_18 ( .A(ab_17__18_), .B(CARRYB_16__18_), .CI(SUMB_16__19_), .CO(
        CARRYB_17__18_), .S(SUMB_17__18_) );
  FA_X1 S2_17_19 ( .A(ab_17__19_), .B(CARRYB_16__19_), .CI(SUMB_16__20_), .CO(
        CARRYB_17__19_), .S(SUMB_17__19_) );
  FA_X1 S2_17_20 ( .A(ab_17__20_), .B(CARRYB_16__20_), .CI(SUMB_16__21_), .CO(
        CARRYB_17__20_), .S(SUMB_17__20_) );
  FA_X1 S2_17_21 ( .A(ab_17__21_), .B(CARRYB_16__21_), .CI(SUMB_16__22_), .CO(
        CARRYB_17__21_), .S(SUMB_17__21_) );
  FA_X1 S3_17_22 ( .A(ab_17__22_), .B(CARRYB_16__22_), .CI(ab_16__23_), .CO(
        CARRYB_17__22_), .S(SUMB_17__22_) );
  FA_X1 S1_16_0 ( .A(ab_16__0_), .B(CARRYB_15__0_), .CI(SUMB_15__1_), .CO(
        CARRYB_16__0_), .S(A1_14_) );
  FA_X1 S2_16_1 ( .A(ab_16__1_), .B(CARRYB_15__1_), .CI(SUMB_15__2_), .CO(
        CARRYB_16__1_), .S(SUMB_16__1_) );
  FA_X1 S2_16_2 ( .A(ab_16__2_), .B(CARRYB_15__2_), .CI(SUMB_15__3_), .CO(
        CARRYB_16__2_), .S(SUMB_16__2_) );
  FA_X1 S2_16_3 ( .A(ab_16__3_), .B(CARRYB_15__3_), .CI(SUMB_15__4_), .CO(
        CARRYB_16__3_), .S(SUMB_16__3_) );
  FA_X1 S2_16_4 ( .A(ab_16__4_), .B(CARRYB_15__4_), .CI(SUMB_15__5_), .CO(
        CARRYB_16__4_), .S(SUMB_16__4_) );
  FA_X1 S2_16_5 ( .A(ab_16__5_), .B(CARRYB_15__5_), .CI(SUMB_15__6_), .CO(
        CARRYB_16__5_), .S(SUMB_16__5_) );
  FA_X1 S2_16_6 ( .A(ab_16__6_), .B(CARRYB_15__6_), .CI(SUMB_15__7_), .CO(
        CARRYB_16__6_), .S(SUMB_16__6_) );
  FA_X1 S2_16_7 ( .A(ab_16__7_), .B(CARRYB_15__7_), .CI(SUMB_15__8_), .CO(
        CARRYB_16__7_), .S(SUMB_16__7_) );
  FA_X1 S2_16_8 ( .A(ab_16__8_), .B(CARRYB_15__8_), .CI(SUMB_15__9_), .CO(
        CARRYB_16__8_), .S(SUMB_16__8_) );
  FA_X1 S2_16_9 ( .A(ab_16__9_), .B(CARRYB_15__9_), .CI(SUMB_15__10_), .CO(
        CARRYB_16__9_), .S(SUMB_16__9_) );
  FA_X1 S2_16_10 ( .A(ab_16__10_), .B(CARRYB_15__10_), .CI(SUMB_15__11_), .CO(
        CARRYB_16__10_), .S(SUMB_16__10_) );
  FA_X1 S2_16_11 ( .A(ab_16__11_), .B(CARRYB_15__11_), .CI(SUMB_15__12_), .CO(
        CARRYB_16__11_), .S(SUMB_16__11_) );
  FA_X1 S2_16_12 ( .A(ab_16__12_), .B(CARRYB_15__12_), .CI(SUMB_15__13_), .CO(
        CARRYB_16__12_), .S(SUMB_16__12_) );
  FA_X1 S2_16_13 ( .A(ab_16__13_), .B(CARRYB_15__13_), .CI(SUMB_15__14_), .CO(
        CARRYB_16__13_), .S(SUMB_16__13_) );
  FA_X1 S2_16_14 ( .A(ab_16__14_), .B(CARRYB_15__14_), .CI(SUMB_15__15_), .CO(
        CARRYB_16__14_), .S(SUMB_16__14_) );
  FA_X1 S2_16_15 ( .A(ab_16__15_), .B(CARRYB_15__15_), .CI(SUMB_15__16_), .CO(
        CARRYB_16__15_), .S(SUMB_16__15_) );
  FA_X1 S2_16_16 ( .A(ab_16__16_), .B(CARRYB_15__16_), .CI(SUMB_15__17_), .CO(
        CARRYB_16__16_), .S(SUMB_16__16_) );
  FA_X1 S2_16_17 ( .A(ab_16__17_), .B(CARRYB_15__17_), .CI(SUMB_15__18_), .CO(
        CARRYB_16__17_), .S(SUMB_16__17_) );
  FA_X1 S2_16_18 ( .A(ab_16__18_), .B(CARRYB_15__18_), .CI(SUMB_15__19_), .CO(
        CARRYB_16__18_), .S(SUMB_16__18_) );
  FA_X1 S2_16_19 ( .A(ab_16__19_), .B(CARRYB_15__19_), .CI(SUMB_15__20_), .CO(
        CARRYB_16__19_), .S(SUMB_16__19_) );
  FA_X1 S2_16_20 ( .A(ab_16__20_), .B(CARRYB_15__20_), .CI(SUMB_15__21_), .CO(
        CARRYB_16__20_), .S(SUMB_16__20_) );
  FA_X1 S2_16_21 ( .A(ab_16__21_), .B(CARRYB_15__21_), .CI(SUMB_15__22_), .CO(
        CARRYB_16__21_), .S(SUMB_16__21_) );
  FA_X1 S3_16_22 ( .A(ab_16__22_), .B(CARRYB_15__22_), .CI(ab_15__23_), .CO(
        CARRYB_16__22_), .S(SUMB_16__22_) );
  FA_X1 S1_15_0 ( .A(ab_15__0_), .B(CARRYB_14__0_), .CI(SUMB_14__1_), .CO(
        CARRYB_15__0_), .S(A1_13_) );
  FA_X1 S2_15_1 ( .A(ab_15__1_), .B(CARRYB_14__1_), .CI(SUMB_14__2_), .CO(
        CARRYB_15__1_), .S(SUMB_15__1_) );
  FA_X1 S2_15_2 ( .A(ab_15__2_), .B(CARRYB_14__2_), .CI(SUMB_14__3_), .CO(
        CARRYB_15__2_), .S(SUMB_15__2_) );
  FA_X1 S2_15_3 ( .A(ab_15__3_), .B(CARRYB_14__3_), .CI(SUMB_14__4_), .CO(
        CARRYB_15__3_), .S(SUMB_15__3_) );
  FA_X1 S2_15_4 ( .A(ab_15__4_), .B(CARRYB_14__4_), .CI(SUMB_14__5_), .CO(
        CARRYB_15__4_), .S(SUMB_15__4_) );
  FA_X1 S2_15_5 ( .A(ab_15__5_), .B(CARRYB_14__5_), .CI(SUMB_14__6_), .CO(
        CARRYB_15__5_), .S(SUMB_15__5_) );
  FA_X1 S2_15_6 ( .A(ab_15__6_), .B(CARRYB_14__6_), .CI(SUMB_14__7_), .CO(
        CARRYB_15__6_), .S(SUMB_15__6_) );
  FA_X1 S2_15_7 ( .A(ab_15__7_), .B(CARRYB_14__7_), .CI(SUMB_14__8_), .CO(
        CARRYB_15__7_), .S(SUMB_15__7_) );
  FA_X1 S2_15_8 ( .A(ab_15__8_), .B(CARRYB_14__8_), .CI(SUMB_14__9_), .CO(
        CARRYB_15__8_), .S(SUMB_15__8_) );
  FA_X1 S2_15_9 ( .A(ab_15__9_), .B(CARRYB_14__9_), .CI(SUMB_14__10_), .CO(
        CARRYB_15__9_), .S(SUMB_15__9_) );
  FA_X1 S2_15_10 ( .A(ab_15__10_), .B(CARRYB_14__10_), .CI(SUMB_14__11_), .CO(
        CARRYB_15__10_), .S(SUMB_15__10_) );
  FA_X1 S2_15_11 ( .A(ab_15__11_), .B(CARRYB_14__11_), .CI(SUMB_14__12_), .CO(
        CARRYB_15__11_), .S(SUMB_15__11_) );
  FA_X1 S2_15_12 ( .A(ab_15__12_), .B(CARRYB_14__12_), .CI(SUMB_14__13_), .CO(
        CARRYB_15__12_), .S(SUMB_15__12_) );
  FA_X1 S2_15_13 ( .A(ab_15__13_), .B(CARRYB_14__13_), .CI(SUMB_14__14_), .CO(
        CARRYB_15__13_), .S(SUMB_15__13_) );
  FA_X1 S2_15_14 ( .A(ab_15__14_), .B(CARRYB_14__14_), .CI(SUMB_14__15_), .CO(
        CARRYB_15__14_), .S(SUMB_15__14_) );
  FA_X1 S2_15_15 ( .A(ab_15__15_), .B(CARRYB_14__15_), .CI(SUMB_14__16_), .CO(
        CARRYB_15__15_), .S(SUMB_15__15_) );
  FA_X1 S2_15_16 ( .A(ab_15__16_), .B(CARRYB_14__16_), .CI(SUMB_14__17_), .CO(
        CARRYB_15__16_), .S(SUMB_15__16_) );
  FA_X1 S2_15_17 ( .A(ab_15__17_), .B(CARRYB_14__17_), .CI(SUMB_14__18_), .CO(
        CARRYB_15__17_), .S(SUMB_15__17_) );
  FA_X1 S2_15_18 ( .A(ab_15__18_), .B(CARRYB_14__18_), .CI(SUMB_14__19_), .CO(
        CARRYB_15__18_), .S(SUMB_15__18_) );
  FA_X1 S2_15_19 ( .A(ab_15__19_), .B(CARRYB_14__19_), .CI(SUMB_14__20_), .CO(
        CARRYB_15__19_), .S(SUMB_15__19_) );
  FA_X1 S2_15_20 ( .A(ab_15__20_), .B(CARRYB_14__20_), .CI(SUMB_14__21_), .CO(
        CARRYB_15__20_), .S(SUMB_15__20_) );
  FA_X1 S2_15_21 ( .A(ab_15__21_), .B(CARRYB_14__21_), .CI(SUMB_14__22_), .CO(
        CARRYB_15__21_), .S(SUMB_15__21_) );
  FA_X1 S3_15_22 ( .A(ab_15__22_), .B(CARRYB_14__22_), .CI(ab_14__23_), .CO(
        CARRYB_15__22_), .S(SUMB_15__22_) );
  FA_X1 S1_14_0 ( .A(ab_14__0_), .B(CARRYB_13__0_), .CI(SUMB_13__1_), .CO(
        CARRYB_14__0_), .S(A1_12_) );
  FA_X1 S2_14_1 ( .A(ab_14__1_), .B(CARRYB_13__1_), .CI(SUMB_13__2_), .CO(
        CARRYB_14__1_), .S(SUMB_14__1_) );
  FA_X1 S2_14_2 ( .A(ab_14__2_), .B(CARRYB_13__2_), .CI(SUMB_13__3_), .CO(
        CARRYB_14__2_), .S(SUMB_14__2_) );
  FA_X1 S2_14_3 ( .A(ab_14__3_), .B(CARRYB_13__3_), .CI(SUMB_13__4_), .CO(
        CARRYB_14__3_), .S(SUMB_14__3_) );
  FA_X1 S2_14_4 ( .A(ab_14__4_), .B(CARRYB_13__4_), .CI(SUMB_13__5_), .CO(
        CARRYB_14__4_), .S(SUMB_14__4_) );
  FA_X1 S2_14_5 ( .A(ab_14__5_), .B(CARRYB_13__5_), .CI(SUMB_13__6_), .CO(
        CARRYB_14__5_), .S(SUMB_14__5_) );
  FA_X1 S2_14_6 ( .A(ab_14__6_), .B(CARRYB_13__6_), .CI(SUMB_13__7_), .CO(
        CARRYB_14__6_), .S(SUMB_14__6_) );
  FA_X1 S2_14_7 ( .A(ab_14__7_), .B(CARRYB_13__7_), .CI(SUMB_13__8_), .CO(
        CARRYB_14__7_), .S(SUMB_14__7_) );
  FA_X1 S2_14_8 ( .A(ab_14__8_), .B(CARRYB_13__8_), .CI(SUMB_13__9_), .CO(
        CARRYB_14__8_), .S(SUMB_14__8_) );
  FA_X1 S2_14_9 ( .A(ab_14__9_), .B(CARRYB_13__9_), .CI(SUMB_13__10_), .CO(
        CARRYB_14__9_), .S(SUMB_14__9_) );
  FA_X1 S2_14_10 ( .A(ab_14__10_), .B(CARRYB_13__10_), .CI(SUMB_13__11_), .CO(
        CARRYB_14__10_), .S(SUMB_14__10_) );
  FA_X1 S2_14_11 ( .A(ab_14__11_), .B(CARRYB_13__11_), .CI(SUMB_13__12_), .CO(
        CARRYB_14__11_), .S(SUMB_14__11_) );
  FA_X1 S2_14_12 ( .A(ab_14__12_), .B(CARRYB_13__12_), .CI(SUMB_13__13_), .CO(
        CARRYB_14__12_), .S(SUMB_14__12_) );
  FA_X1 S2_14_13 ( .A(ab_14__13_), .B(CARRYB_13__13_), .CI(SUMB_13__14_), .CO(
        CARRYB_14__13_), .S(SUMB_14__13_) );
  FA_X1 S2_14_14 ( .A(ab_14__14_), .B(CARRYB_13__14_), .CI(SUMB_13__15_), .CO(
        CARRYB_14__14_), .S(SUMB_14__14_) );
  FA_X1 S2_14_15 ( .A(ab_14__15_), .B(CARRYB_13__15_), .CI(SUMB_13__16_), .CO(
        CARRYB_14__15_), .S(SUMB_14__15_) );
  FA_X1 S2_14_16 ( .A(ab_14__16_), .B(CARRYB_13__16_), .CI(SUMB_13__17_), .CO(
        CARRYB_14__16_), .S(SUMB_14__16_) );
  FA_X1 S2_14_17 ( .A(ab_14__17_), .B(CARRYB_13__17_), .CI(SUMB_13__18_), .CO(
        CARRYB_14__17_), .S(SUMB_14__17_) );
  FA_X1 S2_14_18 ( .A(ab_14__18_), .B(CARRYB_13__18_), .CI(SUMB_13__19_), .CO(
        CARRYB_14__18_), .S(SUMB_14__18_) );
  FA_X1 S2_14_19 ( .A(ab_14__19_), .B(CARRYB_13__19_), .CI(SUMB_13__20_), .CO(
        CARRYB_14__19_), .S(SUMB_14__19_) );
  FA_X1 S2_14_20 ( .A(ab_14__20_), .B(CARRYB_13__20_), .CI(SUMB_13__21_), .CO(
        CARRYB_14__20_), .S(SUMB_14__20_) );
  FA_X1 S2_14_21 ( .A(ab_14__21_), .B(CARRYB_13__21_), .CI(SUMB_13__22_), .CO(
        CARRYB_14__21_), .S(SUMB_14__21_) );
  FA_X1 S3_14_22 ( .A(ab_14__22_), .B(CARRYB_13__22_), .CI(ab_13__23_), .CO(
        CARRYB_14__22_), .S(SUMB_14__22_) );
  FA_X1 S1_13_0 ( .A(ab_13__0_), .B(CARRYB_12__0_), .CI(SUMB_12__1_), .CO(
        CARRYB_13__0_), .S(A1_11_) );
  FA_X1 S2_13_1 ( .A(ab_13__1_), .B(CARRYB_12__1_), .CI(SUMB_12__2_), .CO(
        CARRYB_13__1_), .S(SUMB_13__1_) );
  FA_X1 S2_13_2 ( .A(ab_13__2_), .B(CARRYB_12__2_), .CI(SUMB_12__3_), .CO(
        CARRYB_13__2_), .S(SUMB_13__2_) );
  FA_X1 S2_13_3 ( .A(ab_13__3_), .B(CARRYB_12__3_), .CI(SUMB_12__4_), .CO(
        CARRYB_13__3_), .S(SUMB_13__3_) );
  FA_X1 S2_13_4 ( .A(ab_13__4_), .B(CARRYB_12__4_), .CI(SUMB_12__5_), .CO(
        CARRYB_13__4_), .S(SUMB_13__4_) );
  FA_X1 S2_13_5 ( .A(ab_13__5_), .B(CARRYB_12__5_), .CI(SUMB_12__6_), .CO(
        CARRYB_13__5_), .S(SUMB_13__5_) );
  FA_X1 S2_13_6 ( .A(ab_13__6_), .B(CARRYB_12__6_), .CI(SUMB_12__7_), .CO(
        CARRYB_13__6_), .S(SUMB_13__6_) );
  FA_X1 S2_13_7 ( .A(ab_13__7_), .B(CARRYB_12__7_), .CI(SUMB_12__8_), .CO(
        CARRYB_13__7_), .S(SUMB_13__7_) );
  FA_X1 S2_13_8 ( .A(ab_13__8_), .B(CARRYB_12__8_), .CI(SUMB_12__9_), .CO(
        CARRYB_13__8_), .S(SUMB_13__8_) );
  FA_X1 S2_13_9 ( .A(ab_13__9_), .B(CARRYB_12__9_), .CI(SUMB_12__10_), .CO(
        CARRYB_13__9_), .S(SUMB_13__9_) );
  FA_X1 S2_13_10 ( .A(ab_13__10_), .B(CARRYB_12__10_), .CI(SUMB_12__11_), .CO(
        CARRYB_13__10_), .S(SUMB_13__10_) );
  FA_X1 S2_13_11 ( .A(ab_13__11_), .B(CARRYB_12__11_), .CI(SUMB_12__12_), .CO(
        CARRYB_13__11_), .S(SUMB_13__11_) );
  FA_X1 S2_13_12 ( .A(ab_13__12_), .B(CARRYB_12__12_), .CI(SUMB_12__13_), .CO(
        CARRYB_13__12_), .S(SUMB_13__12_) );
  FA_X1 S2_13_13 ( .A(ab_13__13_), .B(CARRYB_12__13_), .CI(SUMB_12__14_), .CO(
        CARRYB_13__13_), .S(SUMB_13__13_) );
  FA_X1 S2_13_14 ( .A(ab_13__14_), .B(CARRYB_12__14_), .CI(SUMB_12__15_), .CO(
        CARRYB_13__14_), .S(SUMB_13__14_) );
  FA_X1 S2_13_15 ( .A(ab_13__15_), .B(CARRYB_12__15_), .CI(SUMB_12__16_), .CO(
        CARRYB_13__15_), .S(SUMB_13__15_) );
  FA_X1 S2_13_16 ( .A(ab_13__16_), .B(CARRYB_12__16_), .CI(SUMB_12__17_), .CO(
        CARRYB_13__16_), .S(SUMB_13__16_) );
  FA_X1 S2_13_17 ( .A(ab_13__17_), .B(CARRYB_12__17_), .CI(SUMB_12__18_), .CO(
        CARRYB_13__17_), .S(SUMB_13__17_) );
  FA_X1 S2_13_18 ( .A(ab_13__18_), .B(CARRYB_12__18_), .CI(SUMB_12__19_), .CO(
        CARRYB_13__18_), .S(SUMB_13__18_) );
  FA_X1 S2_13_19 ( .A(ab_13__19_), .B(CARRYB_12__19_), .CI(SUMB_12__20_), .CO(
        CARRYB_13__19_), .S(SUMB_13__19_) );
  FA_X1 S2_13_20 ( .A(ab_13__20_), .B(CARRYB_12__20_), .CI(SUMB_12__21_), .CO(
        CARRYB_13__20_), .S(SUMB_13__20_) );
  FA_X1 S2_13_21 ( .A(ab_13__21_), .B(CARRYB_12__21_), .CI(SUMB_12__22_), .CO(
        CARRYB_13__21_), .S(SUMB_13__21_) );
  FA_X1 S3_13_22 ( .A(ab_13__22_), .B(CARRYB_12__22_), .CI(ab_12__23_), .CO(
        CARRYB_13__22_), .S(SUMB_13__22_) );
  FA_X1 S1_12_0 ( .A(ab_12__0_), .B(CARRYB_11__0_), .CI(SUMB_11__1_), .CO(
        CARRYB_12__0_), .S(A1_10_) );
  FA_X1 S2_12_1 ( .A(ab_12__1_), .B(CARRYB_11__1_), .CI(SUMB_11__2_), .CO(
        CARRYB_12__1_), .S(SUMB_12__1_) );
  FA_X1 S2_12_2 ( .A(ab_12__2_), .B(CARRYB_11__2_), .CI(SUMB_11__3_), .CO(
        CARRYB_12__2_), .S(SUMB_12__2_) );
  FA_X1 S2_12_3 ( .A(ab_12__3_), .B(CARRYB_11__3_), .CI(SUMB_11__4_), .CO(
        CARRYB_12__3_), .S(SUMB_12__3_) );
  FA_X1 S2_12_4 ( .A(ab_12__4_), .B(CARRYB_11__4_), .CI(SUMB_11__5_), .CO(
        CARRYB_12__4_), .S(SUMB_12__4_) );
  FA_X1 S2_12_5 ( .A(ab_12__5_), .B(CARRYB_11__5_), .CI(SUMB_11__6_), .CO(
        CARRYB_12__5_), .S(SUMB_12__5_) );
  FA_X1 S2_12_6 ( .A(ab_12__6_), .B(CARRYB_11__6_), .CI(SUMB_11__7_), .CO(
        CARRYB_12__6_), .S(SUMB_12__6_) );
  FA_X1 S2_12_7 ( .A(ab_12__7_), .B(CARRYB_11__7_), .CI(SUMB_11__8_), .CO(
        CARRYB_12__7_), .S(SUMB_12__7_) );
  FA_X1 S2_12_8 ( .A(ab_12__8_), .B(CARRYB_11__8_), .CI(SUMB_11__9_), .CO(
        CARRYB_12__8_), .S(SUMB_12__8_) );
  FA_X1 S2_12_9 ( .A(ab_12__9_), .B(CARRYB_11__9_), .CI(SUMB_11__10_), .CO(
        CARRYB_12__9_), .S(SUMB_12__9_) );
  FA_X1 S2_12_10 ( .A(ab_12__10_), .B(CARRYB_11__10_), .CI(SUMB_11__11_), .CO(
        CARRYB_12__10_), .S(SUMB_12__10_) );
  FA_X1 S2_12_11 ( .A(ab_12__11_), .B(CARRYB_11__11_), .CI(SUMB_11__12_), .CO(
        CARRYB_12__11_), .S(SUMB_12__11_) );
  FA_X1 S2_12_12 ( .A(ab_12__12_), .B(CARRYB_11__12_), .CI(SUMB_11__13_), .CO(
        CARRYB_12__12_), .S(SUMB_12__12_) );
  FA_X1 S2_12_13 ( .A(ab_12__13_), .B(CARRYB_11__13_), .CI(SUMB_11__14_), .CO(
        CARRYB_12__13_), .S(SUMB_12__13_) );
  FA_X1 S2_12_14 ( .A(ab_12__14_), .B(CARRYB_11__14_), .CI(SUMB_11__15_), .CO(
        CARRYB_12__14_), .S(SUMB_12__14_) );
  FA_X1 S2_12_15 ( .A(ab_12__15_), .B(CARRYB_11__15_), .CI(SUMB_11__16_), .CO(
        CARRYB_12__15_), .S(SUMB_12__15_) );
  FA_X1 S2_12_16 ( .A(ab_12__16_), .B(CARRYB_11__16_), .CI(SUMB_11__17_), .CO(
        CARRYB_12__16_), .S(SUMB_12__16_) );
  FA_X1 S2_12_17 ( .A(ab_12__17_), .B(CARRYB_11__17_), .CI(SUMB_11__18_), .CO(
        CARRYB_12__17_), .S(SUMB_12__17_) );
  FA_X1 S2_12_18 ( .A(ab_12__18_), .B(CARRYB_11__18_), .CI(SUMB_11__19_), .CO(
        CARRYB_12__18_), .S(SUMB_12__18_) );
  FA_X1 S2_12_19 ( .A(ab_12__19_), .B(CARRYB_11__19_), .CI(SUMB_11__20_), .CO(
        CARRYB_12__19_), .S(SUMB_12__19_) );
  FA_X1 S2_12_20 ( .A(ab_12__20_), .B(CARRYB_11__20_), .CI(SUMB_11__21_), .CO(
        CARRYB_12__20_), .S(SUMB_12__20_) );
  FA_X1 S2_12_21 ( .A(ab_12__21_), .B(CARRYB_11__21_), .CI(SUMB_11__22_), .CO(
        CARRYB_12__21_), .S(SUMB_12__21_) );
  FA_X1 S3_12_22 ( .A(ab_12__22_), .B(CARRYB_11__22_), .CI(ab_11__23_), .CO(
        CARRYB_12__22_), .S(SUMB_12__22_) );
  FA_X1 S1_11_0 ( .A(ab_11__0_), .B(CARRYB_10__0_), .CI(SUMB_10__1_), .CO(
        CARRYB_11__0_), .S(A1_9_) );
  FA_X1 S2_11_1 ( .A(ab_11__1_), .B(CARRYB_10__1_), .CI(SUMB_10__2_), .CO(
        CARRYB_11__1_), .S(SUMB_11__1_) );
  FA_X1 S2_11_2 ( .A(ab_11__2_), .B(CARRYB_10__2_), .CI(SUMB_10__3_), .CO(
        CARRYB_11__2_), .S(SUMB_11__2_) );
  FA_X1 S2_11_3 ( .A(ab_11__3_), .B(CARRYB_10__3_), .CI(SUMB_10__4_), .CO(
        CARRYB_11__3_), .S(SUMB_11__3_) );
  FA_X1 S2_11_4 ( .A(ab_11__4_), .B(CARRYB_10__4_), .CI(SUMB_10__5_), .CO(
        CARRYB_11__4_), .S(SUMB_11__4_) );
  FA_X1 S2_11_5 ( .A(ab_11__5_), .B(CARRYB_10__5_), .CI(SUMB_10__6_), .CO(
        CARRYB_11__5_), .S(SUMB_11__5_) );
  FA_X1 S2_11_6 ( .A(ab_11__6_), .B(CARRYB_10__6_), .CI(SUMB_10__7_), .CO(
        CARRYB_11__6_), .S(SUMB_11__6_) );
  FA_X1 S2_11_7 ( .A(ab_11__7_), .B(CARRYB_10__7_), .CI(SUMB_10__8_), .CO(
        CARRYB_11__7_), .S(SUMB_11__7_) );
  FA_X1 S2_11_8 ( .A(ab_11__8_), .B(CARRYB_10__8_), .CI(SUMB_10__9_), .CO(
        CARRYB_11__8_), .S(SUMB_11__8_) );
  FA_X1 S2_11_9 ( .A(ab_11__9_), .B(CARRYB_10__9_), .CI(SUMB_10__10_), .CO(
        CARRYB_11__9_), .S(SUMB_11__9_) );
  FA_X1 S2_11_10 ( .A(ab_11__10_), .B(CARRYB_10__10_), .CI(SUMB_10__11_), .CO(
        CARRYB_11__10_), .S(SUMB_11__10_) );
  FA_X1 S2_11_11 ( .A(ab_11__11_), .B(CARRYB_10__11_), .CI(SUMB_10__12_), .CO(
        CARRYB_11__11_), .S(SUMB_11__11_) );
  FA_X1 S2_11_12 ( .A(ab_11__12_), .B(CARRYB_10__12_), .CI(SUMB_10__13_), .CO(
        CARRYB_11__12_), .S(SUMB_11__12_) );
  FA_X1 S2_11_13 ( .A(ab_11__13_), .B(CARRYB_10__13_), .CI(SUMB_10__14_), .CO(
        CARRYB_11__13_), .S(SUMB_11__13_) );
  FA_X1 S2_11_14 ( .A(ab_11__14_), .B(CARRYB_10__14_), .CI(SUMB_10__15_), .CO(
        CARRYB_11__14_), .S(SUMB_11__14_) );
  FA_X1 S2_11_15 ( .A(ab_11__15_), .B(CARRYB_10__15_), .CI(SUMB_10__16_), .CO(
        CARRYB_11__15_), .S(SUMB_11__15_) );
  FA_X1 S2_11_16 ( .A(ab_11__16_), .B(CARRYB_10__16_), .CI(SUMB_10__17_), .CO(
        CARRYB_11__16_), .S(SUMB_11__16_) );
  FA_X1 S2_11_17 ( .A(ab_11__17_), .B(CARRYB_10__17_), .CI(SUMB_10__18_), .CO(
        CARRYB_11__17_), .S(SUMB_11__17_) );
  FA_X1 S2_11_18 ( .A(ab_11__18_), .B(CARRYB_10__18_), .CI(SUMB_10__19_), .CO(
        CARRYB_11__18_), .S(SUMB_11__18_) );
  FA_X1 S2_11_19 ( .A(ab_11__19_), .B(CARRYB_10__19_), .CI(SUMB_10__20_), .CO(
        CARRYB_11__19_), .S(SUMB_11__19_) );
  FA_X1 S2_11_20 ( .A(ab_11__20_), .B(CARRYB_10__20_), .CI(SUMB_10__21_), .CO(
        CARRYB_11__20_), .S(SUMB_11__20_) );
  FA_X1 S2_11_21 ( .A(ab_11__21_), .B(CARRYB_10__21_), .CI(SUMB_10__22_), .CO(
        CARRYB_11__21_), .S(SUMB_11__21_) );
  FA_X1 S3_11_22 ( .A(ab_11__22_), .B(CARRYB_10__22_), .CI(ab_10__23_), .CO(
        CARRYB_11__22_), .S(SUMB_11__22_) );
  FA_X1 S1_10_0 ( .A(ab_10__0_), .B(CARRYB_9__0_), .CI(SUMB_9__1_), .CO(
        CARRYB_10__0_), .S(A1_8_) );
  FA_X1 S2_10_1 ( .A(ab_10__1_), .B(CARRYB_9__1_), .CI(SUMB_9__2_), .CO(
        CARRYB_10__1_), .S(SUMB_10__1_) );
  FA_X1 S2_10_2 ( .A(ab_10__2_), .B(CARRYB_9__2_), .CI(SUMB_9__3_), .CO(
        CARRYB_10__2_), .S(SUMB_10__2_) );
  FA_X1 S2_10_3 ( .A(ab_10__3_), .B(CARRYB_9__3_), .CI(SUMB_9__4_), .CO(
        CARRYB_10__3_), .S(SUMB_10__3_) );
  FA_X1 S2_10_4 ( .A(ab_10__4_), .B(CARRYB_9__4_), .CI(SUMB_9__5_), .CO(
        CARRYB_10__4_), .S(SUMB_10__4_) );
  FA_X1 S2_10_5 ( .A(ab_10__5_), .B(CARRYB_9__5_), .CI(SUMB_9__6_), .CO(
        CARRYB_10__5_), .S(SUMB_10__5_) );
  FA_X1 S2_10_6 ( .A(ab_10__6_), .B(CARRYB_9__6_), .CI(SUMB_9__7_), .CO(
        CARRYB_10__6_), .S(SUMB_10__6_) );
  FA_X1 S2_10_7 ( .A(ab_10__7_), .B(CARRYB_9__7_), .CI(SUMB_9__8_), .CO(
        CARRYB_10__7_), .S(SUMB_10__7_) );
  FA_X1 S2_10_8 ( .A(ab_10__8_), .B(CARRYB_9__8_), .CI(SUMB_9__9_), .CO(
        CARRYB_10__8_), .S(SUMB_10__8_) );
  FA_X1 S2_10_9 ( .A(ab_10__9_), .B(CARRYB_9__9_), .CI(SUMB_9__10_), .CO(
        CARRYB_10__9_), .S(SUMB_10__9_) );
  FA_X1 S2_10_10 ( .A(ab_10__10_), .B(CARRYB_9__10_), .CI(SUMB_9__11_), .CO(
        CARRYB_10__10_), .S(SUMB_10__10_) );
  FA_X1 S2_10_11 ( .A(ab_10__11_), .B(CARRYB_9__11_), .CI(SUMB_9__12_), .CO(
        CARRYB_10__11_), .S(SUMB_10__11_) );
  FA_X1 S2_10_12 ( .A(ab_10__12_), .B(CARRYB_9__12_), .CI(SUMB_9__13_), .CO(
        CARRYB_10__12_), .S(SUMB_10__12_) );
  FA_X1 S2_10_13 ( .A(ab_10__13_), .B(CARRYB_9__13_), .CI(SUMB_9__14_), .CO(
        CARRYB_10__13_), .S(SUMB_10__13_) );
  FA_X1 S2_10_14 ( .A(ab_10__14_), .B(CARRYB_9__14_), .CI(SUMB_9__15_), .CO(
        CARRYB_10__14_), .S(SUMB_10__14_) );
  FA_X1 S2_10_15 ( .A(ab_10__15_), .B(CARRYB_9__15_), .CI(SUMB_9__16_), .CO(
        CARRYB_10__15_), .S(SUMB_10__15_) );
  FA_X1 S2_10_16 ( .A(ab_10__16_), .B(CARRYB_9__16_), .CI(SUMB_9__17_), .CO(
        CARRYB_10__16_), .S(SUMB_10__16_) );
  FA_X1 S2_10_17 ( .A(ab_10__17_), .B(CARRYB_9__17_), .CI(SUMB_9__18_), .CO(
        CARRYB_10__17_), .S(SUMB_10__17_) );
  FA_X1 S2_10_18 ( .A(ab_10__18_), .B(CARRYB_9__18_), .CI(SUMB_9__19_), .CO(
        CARRYB_10__18_), .S(SUMB_10__18_) );
  FA_X1 S2_10_19 ( .A(ab_10__19_), .B(CARRYB_9__19_), .CI(SUMB_9__20_), .CO(
        CARRYB_10__19_), .S(SUMB_10__19_) );
  FA_X1 S2_10_20 ( .A(ab_10__20_), .B(CARRYB_9__20_), .CI(SUMB_9__21_), .CO(
        CARRYB_10__20_), .S(SUMB_10__20_) );
  FA_X1 S2_10_21 ( .A(ab_10__21_), .B(CARRYB_9__21_), .CI(SUMB_9__22_), .CO(
        CARRYB_10__21_), .S(SUMB_10__21_) );
  FA_X1 S3_10_22 ( .A(ab_10__22_), .B(CARRYB_9__22_), .CI(ab_9__23_), .CO(
        CARRYB_10__22_), .S(SUMB_10__22_) );
  FA_X1 S1_9_0 ( .A(ab_9__0_), .B(CARRYB_8__0_), .CI(SUMB_8__1_), .CO(
        CARRYB_9__0_), .S(A1_7_) );
  FA_X1 S2_9_1 ( .A(ab_9__1_), .B(CARRYB_8__1_), .CI(SUMB_8__2_), .CO(
        CARRYB_9__1_), .S(SUMB_9__1_) );
  FA_X1 S2_9_2 ( .A(ab_9__2_), .B(CARRYB_8__2_), .CI(SUMB_8__3_), .CO(
        CARRYB_9__2_), .S(SUMB_9__2_) );
  FA_X1 S2_9_3 ( .A(ab_9__3_), .B(CARRYB_8__3_), .CI(SUMB_8__4_), .CO(
        CARRYB_9__3_), .S(SUMB_9__3_) );
  FA_X1 S2_9_4 ( .A(ab_9__4_), .B(CARRYB_8__4_), .CI(SUMB_8__5_), .CO(
        CARRYB_9__4_), .S(SUMB_9__4_) );
  FA_X1 S2_9_5 ( .A(ab_9__5_), .B(CARRYB_8__5_), .CI(SUMB_8__6_), .CO(
        CARRYB_9__5_), .S(SUMB_9__5_) );
  FA_X1 S2_9_6 ( .A(ab_9__6_), .B(CARRYB_8__6_), .CI(SUMB_8__7_), .CO(
        CARRYB_9__6_), .S(SUMB_9__6_) );
  FA_X1 S2_9_7 ( .A(ab_9__7_), .B(CARRYB_8__7_), .CI(SUMB_8__8_), .CO(
        CARRYB_9__7_), .S(SUMB_9__7_) );
  FA_X1 S2_9_8 ( .A(ab_9__8_), .B(CARRYB_8__8_), .CI(SUMB_8__9_), .CO(
        CARRYB_9__8_), .S(SUMB_9__8_) );
  FA_X1 S2_9_9 ( .A(ab_9__9_), .B(CARRYB_8__9_), .CI(SUMB_8__10_), .CO(
        CARRYB_9__9_), .S(SUMB_9__9_) );
  FA_X1 S2_9_10 ( .A(ab_9__10_), .B(CARRYB_8__10_), .CI(SUMB_8__11_), .CO(
        CARRYB_9__10_), .S(SUMB_9__10_) );
  FA_X1 S2_9_11 ( .A(ab_9__11_), .B(CARRYB_8__11_), .CI(SUMB_8__12_), .CO(
        CARRYB_9__11_), .S(SUMB_9__11_) );
  FA_X1 S2_9_12 ( .A(ab_9__12_), .B(CARRYB_8__12_), .CI(SUMB_8__13_), .CO(
        CARRYB_9__12_), .S(SUMB_9__12_) );
  FA_X1 S2_9_13 ( .A(ab_9__13_), .B(CARRYB_8__13_), .CI(SUMB_8__14_), .CO(
        CARRYB_9__13_), .S(SUMB_9__13_) );
  FA_X1 S2_9_14 ( .A(ab_9__14_), .B(CARRYB_8__14_), .CI(SUMB_8__15_), .CO(
        CARRYB_9__14_), .S(SUMB_9__14_) );
  FA_X1 S2_9_15 ( .A(ab_9__15_), .B(CARRYB_8__15_), .CI(SUMB_8__16_), .CO(
        CARRYB_9__15_), .S(SUMB_9__15_) );
  FA_X1 S2_9_16 ( .A(ab_9__16_), .B(CARRYB_8__16_), .CI(SUMB_8__17_), .CO(
        CARRYB_9__16_), .S(SUMB_9__16_) );
  FA_X1 S2_9_17 ( .A(ab_9__17_), .B(CARRYB_8__17_), .CI(SUMB_8__18_), .CO(
        CARRYB_9__17_), .S(SUMB_9__17_) );
  FA_X1 S2_9_18 ( .A(ab_9__18_), .B(CARRYB_8__18_), .CI(SUMB_8__19_), .CO(
        CARRYB_9__18_), .S(SUMB_9__18_) );
  FA_X1 S2_9_19 ( .A(ab_9__19_), .B(CARRYB_8__19_), .CI(SUMB_8__20_), .CO(
        CARRYB_9__19_), .S(SUMB_9__19_) );
  FA_X1 S2_9_20 ( .A(ab_9__20_), .B(CARRYB_8__20_), .CI(SUMB_8__21_), .CO(
        CARRYB_9__20_), .S(SUMB_9__20_) );
  FA_X1 S2_9_21 ( .A(ab_9__21_), .B(CARRYB_8__21_), .CI(SUMB_8__22_), .CO(
        CARRYB_9__21_), .S(SUMB_9__21_) );
  FA_X1 S3_9_22 ( .A(ab_9__22_), .B(CARRYB_8__22_), .CI(ab_8__23_), .CO(
        CARRYB_9__22_), .S(SUMB_9__22_) );
  FA_X1 S1_8_0 ( .A(ab_8__0_), .B(CARRYB_7__0_), .CI(SUMB_7__1_), .CO(
        CARRYB_8__0_), .S(A1_6_) );
  FA_X1 S2_8_1 ( .A(ab_8__1_), .B(CARRYB_7__1_), .CI(SUMB_7__2_), .CO(
        CARRYB_8__1_), .S(SUMB_8__1_) );
  FA_X1 S2_8_2 ( .A(ab_8__2_), .B(CARRYB_7__2_), .CI(SUMB_7__3_), .CO(
        CARRYB_8__2_), .S(SUMB_8__2_) );
  FA_X1 S2_8_3 ( .A(ab_8__3_), .B(CARRYB_7__3_), .CI(SUMB_7__4_), .CO(
        CARRYB_8__3_), .S(SUMB_8__3_) );
  FA_X1 S2_8_4 ( .A(ab_8__4_), .B(CARRYB_7__4_), .CI(SUMB_7__5_), .CO(
        CARRYB_8__4_), .S(SUMB_8__4_) );
  FA_X1 S2_8_5 ( .A(ab_8__5_), .B(CARRYB_7__5_), .CI(SUMB_7__6_), .CO(
        CARRYB_8__5_), .S(SUMB_8__5_) );
  FA_X1 S2_8_6 ( .A(ab_8__6_), .B(CARRYB_7__6_), .CI(SUMB_7__7_), .CO(
        CARRYB_8__6_), .S(SUMB_8__6_) );
  FA_X1 S2_8_7 ( .A(ab_8__7_), .B(CARRYB_7__7_), .CI(SUMB_7__8_), .CO(
        CARRYB_8__7_), .S(SUMB_8__7_) );
  FA_X1 S2_8_8 ( .A(ab_8__8_), .B(CARRYB_7__8_), .CI(SUMB_7__9_), .CO(
        CARRYB_8__8_), .S(SUMB_8__8_) );
  FA_X1 S2_8_9 ( .A(ab_8__9_), .B(CARRYB_7__9_), .CI(SUMB_7__10_), .CO(
        CARRYB_8__9_), .S(SUMB_8__9_) );
  FA_X1 S2_8_10 ( .A(ab_8__10_), .B(CARRYB_7__10_), .CI(SUMB_7__11_), .CO(
        CARRYB_8__10_), .S(SUMB_8__10_) );
  FA_X1 S2_8_11 ( .A(ab_8__11_), .B(CARRYB_7__11_), .CI(SUMB_7__12_), .CO(
        CARRYB_8__11_), .S(SUMB_8__11_) );
  FA_X1 S2_8_12 ( .A(ab_8__12_), .B(CARRYB_7__12_), .CI(SUMB_7__13_), .CO(
        CARRYB_8__12_), .S(SUMB_8__12_) );
  FA_X1 S2_8_13 ( .A(ab_8__13_), .B(CARRYB_7__13_), .CI(SUMB_7__14_), .CO(
        CARRYB_8__13_), .S(SUMB_8__13_) );
  FA_X1 S2_8_14 ( .A(ab_8__14_), .B(CARRYB_7__14_), .CI(SUMB_7__15_), .CO(
        CARRYB_8__14_), .S(SUMB_8__14_) );
  FA_X1 S2_8_15 ( .A(ab_8__15_), .B(CARRYB_7__15_), .CI(SUMB_7__16_), .CO(
        CARRYB_8__15_), .S(SUMB_8__15_) );
  FA_X1 S2_8_16 ( .A(ab_8__16_), .B(CARRYB_7__16_), .CI(SUMB_7__17_), .CO(
        CARRYB_8__16_), .S(SUMB_8__16_) );
  FA_X1 S2_8_17 ( .A(ab_8__17_), .B(CARRYB_7__17_), .CI(SUMB_7__18_), .CO(
        CARRYB_8__17_), .S(SUMB_8__17_) );
  FA_X1 S2_8_18 ( .A(ab_8__18_), .B(CARRYB_7__18_), .CI(SUMB_7__19_), .CO(
        CARRYB_8__18_), .S(SUMB_8__18_) );
  FA_X1 S2_8_19 ( .A(ab_8__19_), .B(CARRYB_7__19_), .CI(SUMB_7__20_), .CO(
        CARRYB_8__19_), .S(SUMB_8__19_) );
  FA_X1 S2_8_20 ( .A(ab_8__20_), .B(CARRYB_7__20_), .CI(SUMB_7__21_), .CO(
        CARRYB_8__20_), .S(SUMB_8__20_) );
  FA_X1 S2_8_21 ( .A(ab_8__21_), .B(CARRYB_7__21_), .CI(SUMB_7__22_), .CO(
        CARRYB_8__21_), .S(SUMB_8__21_) );
  FA_X1 S3_8_22 ( .A(ab_8__22_), .B(CARRYB_7__22_), .CI(ab_7__23_), .CO(
        CARRYB_8__22_), .S(SUMB_8__22_) );
  FA_X1 S1_7_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(A1_5_) );
  FA_X1 S2_7_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S2_7_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S2_7_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S2_7_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S2_7_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S2_7_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(SUMB_6__7_), .CO(
        CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S2_7_7 ( .A(ab_7__7_), .B(CARRYB_6__7_), .CI(SUMB_6__8_), .CO(
        CARRYB_7__7_), .S(SUMB_7__7_) );
  FA_X1 S2_7_8 ( .A(ab_7__8_), .B(CARRYB_6__8_), .CI(SUMB_6__9_), .CO(
        CARRYB_7__8_), .S(SUMB_7__8_) );
  FA_X1 S2_7_9 ( .A(ab_7__9_), .B(CARRYB_6__9_), .CI(SUMB_6__10_), .CO(
        CARRYB_7__9_), .S(SUMB_7__9_) );
  FA_X1 S2_7_10 ( .A(ab_7__10_), .B(CARRYB_6__10_), .CI(SUMB_6__11_), .CO(
        CARRYB_7__10_), .S(SUMB_7__10_) );
  FA_X1 S2_7_11 ( .A(ab_7__11_), .B(CARRYB_6__11_), .CI(SUMB_6__12_), .CO(
        CARRYB_7__11_), .S(SUMB_7__11_) );
  FA_X1 S2_7_12 ( .A(ab_7__12_), .B(CARRYB_6__12_), .CI(SUMB_6__13_), .CO(
        CARRYB_7__12_), .S(SUMB_7__12_) );
  FA_X1 S2_7_13 ( .A(ab_7__13_), .B(CARRYB_6__13_), .CI(SUMB_6__14_), .CO(
        CARRYB_7__13_), .S(SUMB_7__13_) );
  FA_X1 S2_7_14 ( .A(ab_7__14_), .B(CARRYB_6__14_), .CI(SUMB_6__15_), .CO(
        CARRYB_7__14_), .S(SUMB_7__14_) );
  FA_X1 S2_7_15 ( .A(ab_7__15_), .B(CARRYB_6__15_), .CI(SUMB_6__16_), .CO(
        CARRYB_7__15_), .S(SUMB_7__15_) );
  FA_X1 S2_7_16 ( .A(ab_7__16_), .B(CARRYB_6__16_), .CI(SUMB_6__17_), .CO(
        CARRYB_7__16_), .S(SUMB_7__16_) );
  FA_X1 S2_7_17 ( .A(ab_7__17_), .B(CARRYB_6__17_), .CI(SUMB_6__18_), .CO(
        CARRYB_7__17_), .S(SUMB_7__17_) );
  FA_X1 S2_7_18 ( .A(ab_7__18_), .B(CARRYB_6__18_), .CI(SUMB_6__19_), .CO(
        CARRYB_7__18_), .S(SUMB_7__18_) );
  FA_X1 S2_7_19 ( .A(ab_7__19_), .B(CARRYB_6__19_), .CI(SUMB_6__20_), .CO(
        CARRYB_7__19_), .S(SUMB_7__19_) );
  FA_X1 S2_7_20 ( .A(ab_7__20_), .B(CARRYB_6__20_), .CI(SUMB_6__21_), .CO(
        CARRYB_7__20_), .S(SUMB_7__20_) );
  FA_X1 S2_7_21 ( .A(ab_7__21_), .B(CARRYB_6__21_), .CI(SUMB_6__22_), .CO(
        CARRYB_7__21_), .S(SUMB_7__21_) );
  FA_X1 S3_7_22 ( .A(ab_7__22_), .B(CARRYB_6__22_), .CI(ab_6__23_), .CO(
        CARRYB_7__22_), .S(SUMB_7__22_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S2_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(SUMB_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S2_6_7 ( .A(ab_6__7_), .B(CARRYB_5__7_), .CI(SUMB_5__8_), .CO(
        CARRYB_6__7_), .S(SUMB_6__7_) );
  FA_X1 S2_6_8 ( .A(ab_6__8_), .B(CARRYB_5__8_), .CI(SUMB_5__9_), .CO(
        CARRYB_6__8_), .S(SUMB_6__8_) );
  FA_X1 S2_6_9 ( .A(ab_6__9_), .B(CARRYB_5__9_), .CI(SUMB_5__10_), .CO(
        CARRYB_6__9_), .S(SUMB_6__9_) );
  FA_X1 S2_6_10 ( .A(ab_6__10_), .B(CARRYB_5__10_), .CI(SUMB_5__11_), .CO(
        CARRYB_6__10_), .S(SUMB_6__10_) );
  FA_X1 S2_6_11 ( .A(ab_6__11_), .B(CARRYB_5__11_), .CI(SUMB_5__12_), .CO(
        CARRYB_6__11_), .S(SUMB_6__11_) );
  FA_X1 S2_6_12 ( .A(ab_6__12_), .B(CARRYB_5__12_), .CI(SUMB_5__13_), .CO(
        CARRYB_6__12_), .S(SUMB_6__12_) );
  FA_X1 S2_6_13 ( .A(ab_6__13_), .B(CARRYB_5__13_), .CI(SUMB_5__14_), .CO(
        CARRYB_6__13_), .S(SUMB_6__13_) );
  FA_X1 S2_6_14 ( .A(ab_6__14_), .B(CARRYB_5__14_), .CI(SUMB_5__15_), .CO(
        CARRYB_6__14_), .S(SUMB_6__14_) );
  FA_X1 S2_6_15 ( .A(ab_6__15_), .B(CARRYB_5__15_), .CI(SUMB_5__16_), .CO(
        CARRYB_6__15_), .S(SUMB_6__15_) );
  FA_X1 S2_6_16 ( .A(ab_6__16_), .B(CARRYB_5__16_), .CI(SUMB_5__17_), .CO(
        CARRYB_6__16_), .S(SUMB_6__16_) );
  FA_X1 S2_6_17 ( .A(ab_6__17_), .B(CARRYB_5__17_), .CI(SUMB_5__18_), .CO(
        CARRYB_6__17_), .S(SUMB_6__17_) );
  FA_X1 S2_6_18 ( .A(ab_6__18_), .B(CARRYB_5__18_), .CI(SUMB_5__19_), .CO(
        CARRYB_6__18_), .S(SUMB_6__18_) );
  FA_X1 S2_6_19 ( .A(ab_6__19_), .B(CARRYB_5__19_), .CI(SUMB_5__20_), .CO(
        CARRYB_6__19_), .S(SUMB_6__19_) );
  FA_X1 S2_6_20 ( .A(ab_6__20_), .B(CARRYB_5__20_), .CI(SUMB_5__21_), .CO(
        CARRYB_6__20_), .S(SUMB_6__20_) );
  FA_X1 S2_6_21 ( .A(ab_6__21_), .B(CARRYB_5__21_), .CI(SUMB_5__22_), .CO(
        CARRYB_6__21_), .S(SUMB_6__21_) );
  FA_X1 S3_6_22 ( .A(ab_6__22_), .B(CARRYB_5__22_), .CI(ab_5__23_), .CO(
        CARRYB_6__22_), .S(SUMB_6__22_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S2_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(SUMB_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S2_5_7 ( .A(ab_5__7_), .B(CARRYB_4__7_), .CI(SUMB_4__8_), .CO(
        CARRYB_5__7_), .S(SUMB_5__7_) );
  FA_X1 S2_5_8 ( .A(ab_5__8_), .B(CARRYB_4__8_), .CI(SUMB_4__9_), .CO(
        CARRYB_5__8_), .S(SUMB_5__8_) );
  FA_X1 S2_5_9 ( .A(ab_5__9_), .B(CARRYB_4__9_), .CI(SUMB_4__10_), .CO(
        CARRYB_5__9_), .S(SUMB_5__9_) );
  FA_X1 S2_5_10 ( .A(ab_5__10_), .B(CARRYB_4__10_), .CI(SUMB_4__11_), .CO(
        CARRYB_5__10_), .S(SUMB_5__10_) );
  FA_X1 S2_5_11 ( .A(ab_5__11_), .B(CARRYB_4__11_), .CI(SUMB_4__12_), .CO(
        CARRYB_5__11_), .S(SUMB_5__11_) );
  FA_X1 S2_5_12 ( .A(ab_5__12_), .B(CARRYB_4__12_), .CI(SUMB_4__13_), .CO(
        CARRYB_5__12_), .S(SUMB_5__12_) );
  FA_X1 S2_5_13 ( .A(ab_5__13_), .B(CARRYB_4__13_), .CI(SUMB_4__14_), .CO(
        CARRYB_5__13_), .S(SUMB_5__13_) );
  FA_X1 S2_5_14 ( .A(ab_5__14_), .B(CARRYB_4__14_), .CI(SUMB_4__15_), .CO(
        CARRYB_5__14_), .S(SUMB_5__14_) );
  FA_X1 S2_5_15 ( .A(ab_5__15_), .B(CARRYB_4__15_), .CI(SUMB_4__16_), .CO(
        CARRYB_5__15_), .S(SUMB_5__15_) );
  FA_X1 S2_5_16 ( .A(ab_5__16_), .B(CARRYB_4__16_), .CI(SUMB_4__17_), .CO(
        CARRYB_5__16_), .S(SUMB_5__16_) );
  FA_X1 S2_5_17 ( .A(ab_5__17_), .B(CARRYB_4__17_), .CI(SUMB_4__18_), .CO(
        CARRYB_5__17_), .S(SUMB_5__17_) );
  FA_X1 S2_5_18 ( .A(ab_5__18_), .B(CARRYB_4__18_), .CI(SUMB_4__19_), .CO(
        CARRYB_5__18_), .S(SUMB_5__18_) );
  FA_X1 S2_5_19 ( .A(ab_5__19_), .B(CARRYB_4__19_), .CI(SUMB_4__20_), .CO(
        CARRYB_5__19_), .S(SUMB_5__19_) );
  FA_X1 S2_5_20 ( .A(ab_5__20_), .B(CARRYB_4__20_), .CI(SUMB_4__21_), .CO(
        CARRYB_5__20_), .S(SUMB_5__20_) );
  FA_X1 S2_5_21 ( .A(ab_5__21_), .B(CARRYB_4__21_), .CI(SUMB_4__22_), .CO(
        CARRYB_5__21_), .S(SUMB_5__21_) );
  FA_X1 S3_5_22 ( .A(ab_5__22_), .B(CARRYB_4__22_), .CI(ab_4__23_), .CO(
        CARRYB_5__22_), .S(SUMB_5__22_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S2_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(SUMB_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S2_4_7 ( .A(ab_4__7_), .B(CARRYB_3__7_), .CI(SUMB_3__8_), .CO(
        CARRYB_4__7_), .S(SUMB_4__7_) );
  FA_X1 S2_4_8 ( .A(ab_4__8_), .B(CARRYB_3__8_), .CI(SUMB_3__9_), .CO(
        CARRYB_4__8_), .S(SUMB_4__8_) );
  FA_X1 S2_4_9 ( .A(ab_4__9_), .B(CARRYB_3__9_), .CI(SUMB_3__10_), .CO(
        CARRYB_4__9_), .S(SUMB_4__9_) );
  FA_X1 S2_4_10 ( .A(ab_4__10_), .B(CARRYB_3__10_), .CI(SUMB_3__11_), .CO(
        CARRYB_4__10_), .S(SUMB_4__10_) );
  FA_X1 S2_4_11 ( .A(ab_4__11_), .B(CARRYB_3__11_), .CI(SUMB_3__12_), .CO(
        CARRYB_4__11_), .S(SUMB_4__11_) );
  FA_X1 S2_4_12 ( .A(ab_4__12_), .B(CARRYB_3__12_), .CI(SUMB_3__13_), .CO(
        CARRYB_4__12_), .S(SUMB_4__12_) );
  FA_X1 S2_4_13 ( .A(ab_4__13_), .B(CARRYB_3__13_), .CI(SUMB_3__14_), .CO(
        CARRYB_4__13_), .S(SUMB_4__13_) );
  FA_X1 S2_4_14 ( .A(ab_4__14_), .B(CARRYB_3__14_), .CI(SUMB_3__15_), .CO(
        CARRYB_4__14_), .S(SUMB_4__14_) );
  FA_X1 S2_4_15 ( .A(ab_4__15_), .B(CARRYB_3__15_), .CI(SUMB_3__16_), .CO(
        CARRYB_4__15_), .S(SUMB_4__15_) );
  FA_X1 S2_4_16 ( .A(ab_4__16_), .B(CARRYB_3__16_), .CI(SUMB_3__17_), .CO(
        CARRYB_4__16_), .S(SUMB_4__16_) );
  FA_X1 S2_4_17 ( .A(ab_4__17_), .B(CARRYB_3__17_), .CI(SUMB_3__18_), .CO(
        CARRYB_4__17_), .S(SUMB_4__17_) );
  FA_X1 S2_4_18 ( .A(ab_4__18_), .B(CARRYB_3__18_), .CI(SUMB_3__19_), .CO(
        CARRYB_4__18_), .S(SUMB_4__18_) );
  FA_X1 S2_4_19 ( .A(ab_4__19_), .B(CARRYB_3__19_), .CI(SUMB_3__20_), .CO(
        CARRYB_4__19_), .S(SUMB_4__19_) );
  FA_X1 S2_4_20 ( .A(ab_4__20_), .B(CARRYB_3__20_), .CI(SUMB_3__21_), .CO(
        CARRYB_4__20_), .S(SUMB_4__20_) );
  FA_X1 S2_4_21 ( .A(ab_4__21_), .B(CARRYB_3__21_), .CI(SUMB_3__22_), .CO(
        CARRYB_4__21_), .S(SUMB_4__21_) );
  FA_X1 S3_4_22 ( .A(ab_4__22_), .B(CARRYB_3__22_), .CI(ab_3__23_), .CO(
        CARRYB_4__22_), .S(SUMB_4__22_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S2_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(SUMB_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S2_3_7 ( .A(ab_3__7_), .B(CARRYB_2__7_), .CI(SUMB_2__8_), .CO(
        CARRYB_3__7_), .S(SUMB_3__7_) );
  FA_X1 S2_3_8 ( .A(ab_3__8_), .B(CARRYB_2__8_), .CI(SUMB_2__9_), .CO(
        CARRYB_3__8_), .S(SUMB_3__8_) );
  FA_X1 S2_3_9 ( .A(ab_3__9_), .B(CARRYB_2__9_), .CI(SUMB_2__10_), .CO(
        CARRYB_3__9_), .S(SUMB_3__9_) );
  FA_X1 S2_3_10 ( .A(ab_3__10_), .B(CARRYB_2__10_), .CI(SUMB_2__11_), .CO(
        CARRYB_3__10_), .S(SUMB_3__10_) );
  FA_X1 S2_3_11 ( .A(ab_3__11_), .B(CARRYB_2__11_), .CI(SUMB_2__12_), .CO(
        CARRYB_3__11_), .S(SUMB_3__11_) );
  FA_X1 S2_3_12 ( .A(ab_3__12_), .B(CARRYB_2__12_), .CI(SUMB_2__13_), .CO(
        CARRYB_3__12_), .S(SUMB_3__12_) );
  FA_X1 S2_3_13 ( .A(ab_3__13_), .B(CARRYB_2__13_), .CI(SUMB_2__14_), .CO(
        CARRYB_3__13_), .S(SUMB_3__13_) );
  FA_X1 S2_3_14 ( .A(ab_3__14_), .B(CARRYB_2__14_), .CI(SUMB_2__15_), .CO(
        CARRYB_3__14_), .S(SUMB_3__14_) );
  FA_X1 S2_3_15 ( .A(ab_3__15_), .B(CARRYB_2__15_), .CI(SUMB_2__16_), .CO(
        CARRYB_3__15_), .S(SUMB_3__15_) );
  FA_X1 S2_3_16 ( .A(ab_3__16_), .B(CARRYB_2__16_), .CI(SUMB_2__17_), .CO(
        CARRYB_3__16_), .S(SUMB_3__16_) );
  FA_X1 S2_3_17 ( .A(ab_3__17_), .B(CARRYB_2__17_), .CI(SUMB_2__18_), .CO(
        CARRYB_3__17_), .S(SUMB_3__17_) );
  FA_X1 S2_3_18 ( .A(ab_3__18_), .B(CARRYB_2__18_), .CI(SUMB_2__19_), .CO(
        CARRYB_3__18_), .S(SUMB_3__18_) );
  FA_X1 S2_3_19 ( .A(ab_3__19_), .B(CARRYB_2__19_), .CI(SUMB_2__20_), .CO(
        CARRYB_3__19_), .S(SUMB_3__19_) );
  FA_X1 S2_3_20 ( .A(ab_3__20_), .B(CARRYB_2__20_), .CI(SUMB_2__21_), .CO(
        CARRYB_3__20_), .S(SUMB_3__20_) );
  FA_X1 S2_3_21 ( .A(ab_3__21_), .B(CARRYB_2__21_), .CI(SUMB_2__22_), .CO(
        CARRYB_3__21_), .S(SUMB_3__21_) );
  FA_X1 S3_3_22 ( .A(ab_3__22_), .B(CARRYB_2__22_), .CI(ab_2__23_), .CO(
        CARRYB_3__22_), .S(SUMB_3__22_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(n89), .CO(CARRYB_2__0_), 
        .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n23), .CI(n44), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n22), .CI(n43), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n21), .CI(n42), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n20), .CI(n41), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n19), .CI(n40), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S2_2_6 ( .A(ab_2__6_), .B(n18), .CI(n39), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  FA_X1 S2_2_7 ( .A(ab_2__7_), .B(n17), .CI(n38), .CO(CARRYB_2__7_), .S(
        SUMB_2__7_) );
  FA_X1 S2_2_8 ( .A(ab_2__8_), .B(n16), .CI(n37), .CO(CARRYB_2__8_), .S(
        SUMB_2__8_) );
  FA_X1 S2_2_9 ( .A(ab_2__9_), .B(n15), .CI(n36), .CO(CARRYB_2__9_), .S(
        SUMB_2__9_) );
  FA_X1 S2_2_10 ( .A(ab_2__10_), .B(n14), .CI(n35), .CO(CARRYB_2__10_), .S(
        SUMB_2__10_) );
  FA_X1 S2_2_11 ( .A(ab_2__11_), .B(n13), .CI(n34), .CO(CARRYB_2__11_), .S(
        SUMB_2__11_) );
  FA_X1 S2_2_12 ( .A(ab_2__12_), .B(n12), .CI(n33), .CO(CARRYB_2__12_), .S(
        SUMB_2__12_) );
  FA_X1 S2_2_13 ( .A(ab_2__13_), .B(n11), .CI(n32), .CO(CARRYB_2__13_), .S(
        SUMB_2__13_) );
  FA_X1 S2_2_14 ( .A(ab_2__14_), .B(n10), .CI(n31), .CO(CARRYB_2__14_), .S(
        SUMB_2__14_) );
  FA_X1 S2_2_15 ( .A(ab_2__15_), .B(n9), .CI(n30), .CO(CARRYB_2__15_), .S(
        SUMB_2__15_) );
  FA_X1 S2_2_16 ( .A(ab_2__16_), .B(n8), .CI(n29), .CO(CARRYB_2__16_), .S(
        SUMB_2__16_) );
  FA_X1 S2_2_17 ( .A(ab_2__17_), .B(n7), .CI(n28), .CO(CARRYB_2__17_), .S(
        SUMB_2__17_) );
  FA_X1 S2_2_18 ( .A(ab_2__18_), .B(n6), .CI(n27), .CO(CARRYB_2__18_), .S(
        SUMB_2__18_) );
  FA_X1 S2_2_19 ( .A(ab_2__19_), .B(n5), .CI(n26), .CO(CARRYB_2__19_), .S(
        SUMB_2__19_) );
  FA_X1 S2_2_20 ( .A(ab_2__20_), .B(n4), .CI(n25), .CO(CARRYB_2__20_), .S(
        SUMB_2__20_) );
  FA_X1 S2_2_21 ( .A(ab_2__21_), .B(n3), .CI(n45), .CO(CARRYB_2__21_), .S(
        SUMB_2__21_) );
  FA_X1 S3_2_22 ( .A(ab_2__22_), .B(n24), .CI(ab_1__23_), .CO(CARRYB_2__22_), 
        .S(SUMB_2__22_) );
  fpMultiplier_DW01_add_2 FS_1 ( .A({1'b0, n75, n78, n84, n77, n83, n76, n65, 
        n52, n63, n47, n67, n51, n66, n50, n64, n49, n62, n48, n60, n46, n61, 
        n88, n92, SUMB_23__0_, A1_20_, A1_19_, A1_18_, A1_17_, A1_16_, A1_15_, 
        A1_14_, A1_13_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, 
        A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_}), .B({n79, n87, n82, n86, 
        n81, n85, n80, n72, n59, n70, n54, n74, n58, n73, n57, n71, n56, n69, 
        n55, n68, n53, n91, n90, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({PRODUCT[47:23], 
        SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, 
        SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, 
        SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, 
        SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11, 
        SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, 
        SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, 
        SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17, 
        SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19, 
        SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21}) );
  INV_X1 U2 ( .A(A[0]), .ZN(n228) );
  INV_X1 U3 ( .A(A[1]), .ZN(n227) );
  BUF_X1 U4 ( .A(n181), .Z(n93) );
  AND2_X1 U5 ( .A1(ab_0__22_), .A2(ab_1__21_), .ZN(n3) );
  AND2_X1 U6 ( .A1(ab_0__21_), .A2(ab_1__20_), .ZN(n4) );
  AND2_X1 U7 ( .A1(ab_0__20_), .A2(ab_1__19_), .ZN(n5) );
  AND2_X1 U8 ( .A1(ab_0__19_), .A2(ab_1__18_), .ZN(n6) );
  AND2_X1 U9 ( .A1(ab_0__18_), .A2(ab_1__17_), .ZN(n7) );
  AND2_X1 U10 ( .A1(ab_0__17_), .A2(ab_1__16_), .ZN(n8) );
  AND2_X1 U11 ( .A1(ab_0__16_), .A2(ab_1__15_), .ZN(n9) );
  AND2_X1 U12 ( .A1(ab_0__15_), .A2(ab_1__14_), .ZN(n10) );
  AND2_X1 U13 ( .A1(ab_0__14_), .A2(ab_1__13_), .ZN(n11) );
  AND2_X1 U14 ( .A1(ab_0__13_), .A2(ab_1__12_), .ZN(n12) );
  AND2_X1 U15 ( .A1(ab_0__12_), .A2(ab_1__11_), .ZN(n13) );
  AND2_X1 U16 ( .A1(ab_0__11_), .A2(ab_1__10_), .ZN(n14) );
  AND2_X1 U17 ( .A1(ab_0__10_), .A2(ab_1__9_), .ZN(n15) );
  AND2_X1 U18 ( .A1(ab_0__9_), .A2(ab_1__8_), .ZN(n16) );
  AND2_X1 U19 ( .A1(ab_0__8_), .A2(ab_1__7_), .ZN(n17) );
  AND2_X1 U20 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n18) );
  AND2_X1 U21 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n19) );
  AND2_X1 U22 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n20) );
  AND2_X1 U23 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n21) );
  AND2_X1 U24 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n22) );
  AND2_X1 U25 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n23) );
  AND2_X1 U26 ( .A1(ab_0__23_), .A2(ab_1__22_), .ZN(n24) );
  XOR2_X1 U27 ( .A(ab_1__21_), .B(ab_0__22_), .Z(n25) );
  XOR2_X1 U28 ( .A(ab_1__20_), .B(ab_0__21_), .Z(n26) );
  XOR2_X1 U29 ( .A(ab_1__19_), .B(ab_0__20_), .Z(n27) );
  XOR2_X1 U30 ( .A(ab_1__18_), .B(ab_0__19_), .Z(n28) );
  XOR2_X1 U31 ( .A(ab_1__17_), .B(ab_0__18_), .Z(n29) );
  XOR2_X1 U32 ( .A(ab_1__16_), .B(ab_0__17_), .Z(n30) );
  XOR2_X1 U33 ( .A(ab_1__15_), .B(ab_0__16_), .Z(n31) );
  XOR2_X1 U34 ( .A(ab_1__14_), .B(ab_0__15_), .Z(n32) );
  XOR2_X1 U35 ( .A(ab_1__13_), .B(ab_0__14_), .Z(n33) );
  XOR2_X1 U36 ( .A(ab_1__12_), .B(ab_0__13_), .Z(n34) );
  XOR2_X1 U37 ( .A(ab_1__11_), .B(ab_0__12_), .Z(n35) );
  XOR2_X1 U38 ( .A(ab_1__10_), .B(ab_0__11_), .Z(n36) );
  XOR2_X1 U39 ( .A(ab_1__9_), .B(ab_0__10_), .Z(n37) );
  XOR2_X1 U40 ( .A(ab_1__8_), .B(ab_0__9_), .Z(n38) );
  XOR2_X1 U41 ( .A(ab_1__7_), .B(ab_0__8_), .Z(n39) );
  XOR2_X1 U42 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n40) );
  XOR2_X1 U43 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n41) );
  XOR2_X1 U44 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n42) );
  XOR2_X1 U45 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n43) );
  XOR2_X1 U46 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n44) );
  XOR2_X1 U47 ( .A(ab_1__22_), .B(ab_0__23_), .Z(n45) );
  XOR2_X1 U48 ( .A(CARRYB_23__3_), .B(SUMB_23__4_), .Z(n46) );
  XOR2_X1 U49 ( .A(CARRYB_23__13_), .B(SUMB_23__14_), .Z(n47) );
  XOR2_X1 U50 ( .A(CARRYB_23__5_), .B(SUMB_23__6_), .Z(n48) );
  XOR2_X1 U51 ( .A(CARRYB_23__7_), .B(SUMB_23__8_), .Z(n49) );
  XOR2_X1 U52 ( .A(CARRYB_23__9_), .B(SUMB_23__10_), .Z(n50) );
  XOR2_X1 U53 ( .A(CARRYB_23__11_), .B(SUMB_23__12_), .Z(n51) );
  XOR2_X1 U54 ( .A(CARRYB_23__15_), .B(SUMB_23__16_), .Z(n52) );
  AND2_X1 U55 ( .A1(CARRYB_23__2_), .A2(SUMB_23__3_), .ZN(n53) );
  AND2_X1 U56 ( .A1(CARRYB_23__12_), .A2(SUMB_23__13_), .ZN(n54) );
  AND2_X1 U57 ( .A1(CARRYB_23__4_), .A2(SUMB_23__5_), .ZN(n55) );
  AND2_X1 U58 ( .A1(CARRYB_23__6_), .A2(SUMB_23__7_), .ZN(n56) );
  AND2_X1 U59 ( .A1(CARRYB_23__8_), .A2(SUMB_23__9_), .ZN(n57) );
  AND2_X1 U60 ( .A1(CARRYB_23__10_), .A2(SUMB_23__11_), .ZN(n58) );
  AND2_X1 U61 ( .A1(CARRYB_23__14_), .A2(SUMB_23__15_), .ZN(n59) );
  XOR2_X1 U62 ( .A(CARRYB_23__4_), .B(SUMB_23__5_), .Z(n60) );
  XOR2_X1 U63 ( .A(CARRYB_23__2_), .B(SUMB_23__3_), .Z(n61) );
  XOR2_X1 U64 ( .A(CARRYB_23__6_), .B(SUMB_23__7_), .Z(n62) );
  XOR2_X1 U65 ( .A(CARRYB_23__14_), .B(SUMB_23__15_), .Z(n63) );
  XOR2_X1 U66 ( .A(CARRYB_23__8_), .B(SUMB_23__9_), .Z(n64) );
  XOR2_X1 U67 ( .A(CARRYB_23__16_), .B(SUMB_23__17_), .Z(n65) );
  XOR2_X1 U68 ( .A(CARRYB_23__10_), .B(SUMB_23__11_), .Z(n66) );
  XOR2_X1 U69 ( .A(CARRYB_23__12_), .B(SUMB_23__13_), .Z(n67) );
  AND2_X1 U70 ( .A1(CARRYB_23__3_), .A2(SUMB_23__4_), .ZN(n68) );
  AND2_X1 U71 ( .A1(CARRYB_23__5_), .A2(SUMB_23__6_), .ZN(n69) );
  AND2_X1 U72 ( .A1(CARRYB_23__13_), .A2(SUMB_23__14_), .ZN(n70) );
  AND2_X1 U73 ( .A1(CARRYB_23__7_), .A2(SUMB_23__8_), .ZN(n71) );
  AND2_X1 U74 ( .A1(CARRYB_23__15_), .A2(SUMB_23__16_), .ZN(n72) );
  AND2_X1 U75 ( .A1(CARRYB_23__9_), .A2(SUMB_23__10_), .ZN(n73) );
  AND2_X1 U76 ( .A1(CARRYB_23__11_), .A2(SUMB_23__12_), .ZN(n74) );
  XOR2_X1 U77 ( .A(CARRYB_23__22_), .B(ab_23__23_), .Z(n75) );
  XOR2_X1 U78 ( .A(CARRYB_23__17_), .B(SUMB_23__18_), .Z(n76) );
  XOR2_X1 U79 ( .A(CARRYB_23__19_), .B(SUMB_23__20_), .Z(n77) );
  XOR2_X1 U80 ( .A(CARRYB_23__21_), .B(SUMB_23__22_), .Z(n78) );
  AND2_X1 U81 ( .A1(CARRYB_23__22_), .A2(ab_23__23_), .ZN(n79) );
  AND2_X1 U82 ( .A1(CARRYB_23__16_), .A2(SUMB_23__17_), .ZN(n80) );
  AND2_X1 U83 ( .A1(CARRYB_23__18_), .A2(SUMB_23__19_), .ZN(n81) );
  AND2_X1 U84 ( .A1(CARRYB_23__20_), .A2(SUMB_23__21_), .ZN(n82) );
  XOR2_X1 U85 ( .A(CARRYB_23__18_), .B(SUMB_23__19_), .Z(n83) );
  XOR2_X1 U86 ( .A(CARRYB_23__20_), .B(SUMB_23__21_), .Z(n84) );
  AND2_X1 U87 ( .A1(CARRYB_23__17_), .A2(SUMB_23__18_), .ZN(n85) );
  AND2_X1 U88 ( .A1(CARRYB_23__19_), .A2(SUMB_23__20_), .ZN(n86) );
  AND2_X1 U89 ( .A1(CARRYB_23__21_), .A2(SUMB_23__22_), .ZN(n87) );
  BUF_X1 U90 ( .A(n181), .Z(n94) );
  XOR2_X1 U91 ( .A(CARRYB_23__1_), .B(SUMB_23__2_), .Z(n88) );
  XOR2_X1 U92 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n89) );
  AND2_X1 U93 ( .A1(CARRYB_23__0_), .A2(SUMB_23__1_), .ZN(n90) );
  AND2_X1 U94 ( .A1(CARRYB_23__1_), .A2(SUMB_23__2_), .ZN(n91) );
  XOR2_X1 U95 ( .A(CARRYB_23__0_), .B(SUMB_23__1_), .Z(n92) );
  BUF_X1 U96 ( .A(n205), .Z(n137) );
  BUF_X1 U97 ( .A(n205), .Z(n138) );
  BUF_X1 U98 ( .A(n184), .Z(n99) );
  BUF_X1 U99 ( .A(n183), .Z(n97) );
  BUF_X1 U100 ( .A(n182), .Z(n95) );
  BUF_X1 U101 ( .A(n185), .Z(n101) );
  BUF_X1 U102 ( .A(n186), .Z(n103) );
  BUF_X1 U103 ( .A(n187), .Z(n105) );
  BUF_X1 U104 ( .A(n188), .Z(n107) );
  BUF_X1 U105 ( .A(n189), .Z(n109) );
  BUF_X1 U106 ( .A(n190), .Z(n111) );
  BUF_X1 U107 ( .A(n191), .Z(n113) );
  BUF_X1 U108 ( .A(n192), .Z(n115) );
  BUF_X1 U109 ( .A(n193), .Z(n117) );
  BUF_X1 U110 ( .A(n194), .Z(n119) );
  BUF_X1 U111 ( .A(n195), .Z(n121) );
  BUF_X1 U112 ( .A(n196), .Z(n123) );
  BUF_X1 U113 ( .A(n197), .Z(n125) );
  BUF_X1 U114 ( .A(n198), .Z(n127) );
  BUF_X1 U115 ( .A(n199), .Z(n129) );
  BUF_X1 U116 ( .A(n200), .Z(n131) );
  BUF_X1 U117 ( .A(n202), .Z(n135) );
  BUF_X1 U118 ( .A(n201), .Z(n133) );
  BUF_X1 U119 ( .A(n188), .Z(n108) );
  BUF_X1 U120 ( .A(n202), .Z(n136) );
  BUF_X1 U121 ( .A(n189), .Z(n110) );
  BUF_X1 U122 ( .A(n190), .Z(n112) );
  BUF_X1 U123 ( .A(n191), .Z(n114) );
  BUF_X1 U124 ( .A(n192), .Z(n116) );
  BUF_X1 U125 ( .A(n193), .Z(n118) );
  BUF_X1 U126 ( .A(n194), .Z(n120) );
  BUF_X1 U127 ( .A(n195), .Z(n122) );
  BUF_X1 U128 ( .A(n196), .Z(n124) );
  BUF_X1 U129 ( .A(n197), .Z(n126) );
  BUF_X1 U130 ( .A(n198), .Z(n128) );
  BUF_X1 U131 ( .A(n199), .Z(n130) );
  BUF_X1 U132 ( .A(n200), .Z(n132) );
  BUF_X1 U133 ( .A(n201), .Z(n134) );
  BUF_X1 U134 ( .A(n186), .Z(n104) );
  BUF_X1 U135 ( .A(n187), .Z(n106) );
  BUF_X1 U136 ( .A(n185), .Z(n102) );
  BUF_X1 U137 ( .A(n184), .Z(n100) );
  BUF_X1 U138 ( .A(n182), .Z(n96) );
  BUF_X1 U139 ( .A(n183), .Z(n98) );
  BUF_X1 U140 ( .A(n226), .Z(n180) );
  BUF_X1 U141 ( .A(n225), .Z(n178) );
  BUF_X1 U142 ( .A(n224), .Z(n176) );
  BUF_X1 U143 ( .A(n223), .Z(n174) );
  BUF_X1 U144 ( .A(n222), .Z(n172) );
  BUF_X1 U145 ( .A(n221), .Z(n170) );
  BUF_X1 U146 ( .A(n220), .Z(n168) );
  BUF_X1 U147 ( .A(n226), .Z(n179) );
  BUF_X1 U148 ( .A(n225), .Z(n177) );
  BUF_X1 U149 ( .A(n224), .Z(n175) );
  BUF_X1 U150 ( .A(n223), .Z(n173) );
  BUF_X1 U151 ( .A(n222), .Z(n171) );
  BUF_X1 U152 ( .A(n221), .Z(n169) );
  BUF_X1 U153 ( .A(n220), .Z(n167) );
  BUF_X1 U154 ( .A(n219), .Z(n166) );
  BUF_X1 U155 ( .A(n219), .Z(n165) );
  BUF_X1 U156 ( .A(n218), .Z(n164) );
  BUF_X1 U157 ( .A(n217), .Z(n162) );
  BUF_X1 U158 ( .A(n216), .Z(n160) );
  BUF_X1 U159 ( .A(n215), .Z(n158) );
  BUF_X1 U160 ( .A(n214), .Z(n156) );
  BUF_X1 U161 ( .A(n213), .Z(n154) );
  BUF_X1 U162 ( .A(n212), .Z(n152) );
  BUF_X1 U163 ( .A(n211), .Z(n150) );
  BUF_X1 U164 ( .A(n218), .Z(n163) );
  BUF_X1 U165 ( .A(n217), .Z(n161) );
  BUF_X1 U166 ( .A(n216), .Z(n159) );
  BUF_X1 U167 ( .A(n215), .Z(n157) );
  BUF_X1 U168 ( .A(n214), .Z(n155) );
  BUF_X1 U169 ( .A(n213), .Z(n153) );
  BUF_X1 U170 ( .A(n212), .Z(n151) );
  BUF_X1 U171 ( .A(n211), .Z(n149) );
  BUF_X1 U172 ( .A(n210), .Z(n148) );
  BUF_X1 U173 ( .A(n209), .Z(n146) );
  BUF_X1 U174 ( .A(n208), .Z(n144) );
  BUF_X1 U175 ( .A(n207), .Z(n142) );
  BUF_X1 U176 ( .A(n206), .Z(n140) );
  BUF_X1 U177 ( .A(n210), .Z(n147) );
  BUF_X1 U178 ( .A(n209), .Z(n145) );
  BUF_X1 U179 ( .A(n208), .Z(n143) );
  BUF_X1 U180 ( .A(n207), .Z(n141) );
  BUF_X1 U181 ( .A(n206), .Z(n139) );
  INV_X1 U182 ( .A(A[23]), .ZN(n205) );
  INV_X1 U183 ( .A(B[1]), .ZN(n203) );
  INV_X1 U184 ( .A(B[0]), .ZN(n204) );
  INV_X1 U185 ( .A(B[20]), .ZN(n184) );
  INV_X1 U186 ( .A(B[15]), .ZN(n189) );
  INV_X1 U187 ( .A(B[5]), .ZN(n199) );
  INV_X1 U188 ( .A(A[5]), .ZN(n223) );
  INV_X1 U189 ( .A(B[21]), .ZN(n183) );
  INV_X1 U190 ( .A(B[16]), .ZN(n188) );
  INV_X1 U191 ( .A(B[10]), .ZN(n194) );
  INV_X1 U192 ( .A(B[6]), .ZN(n198) );
  INV_X1 U193 ( .A(A[6]), .ZN(n222) );
  INV_X1 U194 ( .A(B[14]), .ZN(n190) );
  INV_X1 U195 ( .A(B[4]), .ZN(n200) );
  INV_X1 U196 ( .A(A[4]), .ZN(n224) );
  INV_X1 U197 ( .A(B[22]), .ZN(n182) );
  INV_X1 U198 ( .A(B[19]), .ZN(n185) );
  INV_X1 U199 ( .A(B[18]), .ZN(n186) );
  INV_X1 U200 ( .A(B[17]), .ZN(n187) );
  INV_X1 U201 ( .A(B[13]), .ZN(n191) );
  INV_X1 U202 ( .A(B[12]), .ZN(n192) );
  INV_X1 U203 ( .A(B[11]), .ZN(n193) );
  INV_X1 U204 ( .A(B[9]), .ZN(n195) );
  INV_X1 U205 ( .A(B[8]), .ZN(n196) );
  INV_X1 U206 ( .A(B[7]), .ZN(n197) );
  INV_X1 U207 ( .A(B[2]), .ZN(n202) );
  INV_X1 U208 ( .A(B[3]), .ZN(n201) );
  INV_X1 U209 ( .A(A[2]), .ZN(n226) );
  INV_X1 U210 ( .A(A[3]), .ZN(n225) );
  INV_X1 U211 ( .A(A[7]), .ZN(n221) );
  INV_X1 U212 ( .A(A[8]), .ZN(n220) );
  INV_X1 U213 ( .A(A[15]), .ZN(n213) );
  INV_X1 U214 ( .A(A[10]), .ZN(n218) );
  INV_X1 U215 ( .A(A[16]), .ZN(n212) );
  INV_X1 U216 ( .A(A[14]), .ZN(n214) );
  INV_X1 U217 ( .A(A[9]), .ZN(n219) );
  INV_X1 U218 ( .A(A[11]), .ZN(n217) );
  INV_X1 U219 ( .A(A[12]), .ZN(n216) );
  INV_X1 U220 ( .A(A[13]), .ZN(n215) );
  INV_X1 U221 ( .A(A[17]), .ZN(n211) );
  INV_X1 U222 ( .A(A[20]), .ZN(n208) );
  INV_X1 U223 ( .A(A[21]), .ZN(n207) );
  INV_X1 U224 ( .A(A[18]), .ZN(n210) );
  INV_X1 U225 ( .A(A[19]), .ZN(n209) );
  INV_X1 U226 ( .A(A[22]), .ZN(n206) );
  INV_X1 U227 ( .A(B[23]), .ZN(n181) );
  NOR2_X1 U229 ( .A1(n166), .A2(n122), .ZN(ab_9__9_) );
  NOR2_X1 U230 ( .A1(n166), .A2(n124), .ZN(ab_9__8_) );
  NOR2_X1 U231 ( .A1(n166), .A2(n126), .ZN(ab_9__7_) );
  NOR2_X1 U232 ( .A1(n166), .A2(n128), .ZN(ab_9__6_) );
  NOR2_X1 U233 ( .A1(n166), .A2(n130), .ZN(ab_9__5_) );
  NOR2_X1 U234 ( .A1(n166), .A2(n132), .ZN(ab_9__4_) );
  NOR2_X1 U235 ( .A1(n166), .A2(n134), .ZN(ab_9__3_) );
  NOR2_X1 U236 ( .A1(n166), .A2(n136), .ZN(ab_9__2_) );
  NOR2_X1 U237 ( .A1(n166), .A2(n94), .ZN(ab_9__23_) );
  NOR2_X1 U238 ( .A1(n166), .A2(n96), .ZN(ab_9__22_) );
  NOR2_X1 U239 ( .A1(n166), .A2(n98), .ZN(ab_9__21_) );
  NOR2_X1 U240 ( .A1(n166), .A2(n100), .ZN(ab_9__20_) );
  NOR2_X1 U241 ( .A1(n165), .A2(n203), .ZN(ab_9__1_) );
  NOR2_X1 U242 ( .A1(n165), .A2(n102), .ZN(ab_9__19_) );
  NOR2_X1 U243 ( .A1(n165), .A2(n104), .ZN(ab_9__18_) );
  NOR2_X1 U244 ( .A1(n165), .A2(n106), .ZN(ab_9__17_) );
  NOR2_X1 U245 ( .A1(n165), .A2(n108), .ZN(ab_9__16_) );
  NOR2_X1 U246 ( .A1(n165), .A2(n110), .ZN(ab_9__15_) );
  NOR2_X1 U247 ( .A1(n165), .A2(n112), .ZN(ab_9__14_) );
  NOR2_X1 U248 ( .A1(n165), .A2(n114), .ZN(ab_9__13_) );
  NOR2_X1 U249 ( .A1(n165), .A2(n116), .ZN(ab_9__12_) );
  NOR2_X1 U250 ( .A1(n165), .A2(n118), .ZN(ab_9__11_) );
  NOR2_X1 U251 ( .A1(n165), .A2(n120), .ZN(ab_9__10_) );
  NOR2_X1 U252 ( .A1(n165), .A2(n204), .ZN(ab_9__0_) );
  NOR2_X1 U253 ( .A1(n122), .A2(n168), .ZN(ab_8__9_) );
  NOR2_X1 U254 ( .A1(n124), .A2(n168), .ZN(ab_8__8_) );
  NOR2_X1 U255 ( .A1(n126), .A2(n168), .ZN(ab_8__7_) );
  NOR2_X1 U256 ( .A1(n128), .A2(n168), .ZN(ab_8__6_) );
  NOR2_X1 U257 ( .A1(n130), .A2(n168), .ZN(ab_8__5_) );
  NOR2_X1 U258 ( .A1(n132), .A2(n168), .ZN(ab_8__4_) );
  NOR2_X1 U259 ( .A1(n134), .A2(n168), .ZN(ab_8__3_) );
  NOR2_X1 U260 ( .A1(n136), .A2(n168), .ZN(ab_8__2_) );
  NOR2_X1 U261 ( .A1(n94), .A2(n168), .ZN(ab_8__23_) );
  NOR2_X1 U262 ( .A1(n96), .A2(n168), .ZN(ab_8__22_) );
  NOR2_X1 U263 ( .A1(n98), .A2(n168), .ZN(ab_8__21_) );
  NOR2_X1 U264 ( .A1(n100), .A2(n168), .ZN(ab_8__20_) );
  NOR2_X1 U265 ( .A1(n203), .A2(n167), .ZN(ab_8__1_) );
  NOR2_X1 U266 ( .A1(n102), .A2(n167), .ZN(ab_8__19_) );
  NOR2_X1 U267 ( .A1(n104), .A2(n167), .ZN(ab_8__18_) );
  NOR2_X1 U268 ( .A1(n106), .A2(n167), .ZN(ab_8__17_) );
  NOR2_X1 U269 ( .A1(n108), .A2(n167), .ZN(ab_8__16_) );
  NOR2_X1 U270 ( .A1(n110), .A2(n167), .ZN(ab_8__15_) );
  NOR2_X1 U271 ( .A1(n112), .A2(n167), .ZN(ab_8__14_) );
  NOR2_X1 U272 ( .A1(n114), .A2(n167), .ZN(ab_8__13_) );
  NOR2_X1 U273 ( .A1(n116), .A2(n167), .ZN(ab_8__12_) );
  NOR2_X1 U274 ( .A1(n118), .A2(n167), .ZN(ab_8__11_) );
  NOR2_X1 U275 ( .A1(n120), .A2(n167), .ZN(ab_8__10_) );
  NOR2_X1 U276 ( .A1(n204), .A2(n167), .ZN(ab_8__0_) );
  NOR2_X1 U277 ( .A1(n122), .A2(n170), .ZN(ab_7__9_) );
  NOR2_X1 U278 ( .A1(n124), .A2(n170), .ZN(ab_7__8_) );
  NOR2_X1 U279 ( .A1(n126), .A2(n170), .ZN(ab_7__7_) );
  NOR2_X1 U280 ( .A1(n128), .A2(n170), .ZN(ab_7__6_) );
  NOR2_X1 U281 ( .A1(n130), .A2(n170), .ZN(ab_7__5_) );
  NOR2_X1 U282 ( .A1(n132), .A2(n170), .ZN(ab_7__4_) );
  NOR2_X1 U283 ( .A1(n134), .A2(n170), .ZN(ab_7__3_) );
  NOR2_X1 U284 ( .A1(n136), .A2(n170), .ZN(ab_7__2_) );
  NOR2_X1 U285 ( .A1(n94), .A2(n170), .ZN(ab_7__23_) );
  NOR2_X1 U286 ( .A1(n96), .A2(n170), .ZN(ab_7__22_) );
  NOR2_X1 U287 ( .A1(n98), .A2(n170), .ZN(ab_7__21_) );
  NOR2_X1 U288 ( .A1(n100), .A2(n170), .ZN(ab_7__20_) );
  NOR2_X1 U289 ( .A1(n203), .A2(n169), .ZN(ab_7__1_) );
  NOR2_X1 U290 ( .A1(n102), .A2(n169), .ZN(ab_7__19_) );
  NOR2_X1 U291 ( .A1(n104), .A2(n169), .ZN(ab_7__18_) );
  NOR2_X1 U292 ( .A1(n106), .A2(n169), .ZN(ab_7__17_) );
  NOR2_X1 U293 ( .A1(n108), .A2(n169), .ZN(ab_7__16_) );
  NOR2_X1 U294 ( .A1(n110), .A2(n169), .ZN(ab_7__15_) );
  NOR2_X1 U295 ( .A1(n112), .A2(n169), .ZN(ab_7__14_) );
  NOR2_X1 U296 ( .A1(n114), .A2(n169), .ZN(ab_7__13_) );
  NOR2_X1 U297 ( .A1(n116), .A2(n169), .ZN(ab_7__12_) );
  NOR2_X1 U298 ( .A1(n118), .A2(n169), .ZN(ab_7__11_) );
  NOR2_X1 U299 ( .A1(n120), .A2(n169), .ZN(ab_7__10_) );
  NOR2_X1 U300 ( .A1(n204), .A2(n169), .ZN(ab_7__0_) );
  NOR2_X1 U301 ( .A1(n122), .A2(n172), .ZN(ab_6__9_) );
  NOR2_X1 U302 ( .A1(n124), .A2(n172), .ZN(ab_6__8_) );
  NOR2_X1 U303 ( .A1(n126), .A2(n172), .ZN(ab_6__7_) );
  NOR2_X1 U304 ( .A1(n128), .A2(n172), .ZN(ab_6__6_) );
  NOR2_X1 U305 ( .A1(n130), .A2(n172), .ZN(ab_6__5_) );
  NOR2_X1 U306 ( .A1(n132), .A2(n172), .ZN(ab_6__4_) );
  NOR2_X1 U307 ( .A1(n134), .A2(n172), .ZN(ab_6__3_) );
  NOR2_X1 U308 ( .A1(n136), .A2(n172), .ZN(ab_6__2_) );
  NOR2_X1 U309 ( .A1(n94), .A2(n172), .ZN(ab_6__23_) );
  NOR2_X1 U310 ( .A1(n96), .A2(n172), .ZN(ab_6__22_) );
  NOR2_X1 U311 ( .A1(n98), .A2(n172), .ZN(ab_6__21_) );
  NOR2_X1 U312 ( .A1(n100), .A2(n172), .ZN(ab_6__20_) );
  NOR2_X1 U313 ( .A1(n203), .A2(n171), .ZN(ab_6__1_) );
  NOR2_X1 U314 ( .A1(n102), .A2(n171), .ZN(ab_6__19_) );
  NOR2_X1 U315 ( .A1(n104), .A2(n171), .ZN(ab_6__18_) );
  NOR2_X1 U316 ( .A1(n106), .A2(n171), .ZN(ab_6__17_) );
  NOR2_X1 U317 ( .A1(n108), .A2(n171), .ZN(ab_6__16_) );
  NOR2_X1 U318 ( .A1(n110), .A2(n171), .ZN(ab_6__15_) );
  NOR2_X1 U319 ( .A1(n112), .A2(n171), .ZN(ab_6__14_) );
  NOR2_X1 U320 ( .A1(n114), .A2(n171), .ZN(ab_6__13_) );
  NOR2_X1 U321 ( .A1(n116), .A2(n171), .ZN(ab_6__12_) );
  NOR2_X1 U322 ( .A1(n118), .A2(n171), .ZN(ab_6__11_) );
  NOR2_X1 U323 ( .A1(n120), .A2(n171), .ZN(ab_6__10_) );
  NOR2_X1 U324 ( .A1(n204), .A2(n171), .ZN(ab_6__0_) );
  NOR2_X1 U325 ( .A1(n122), .A2(n174), .ZN(ab_5__9_) );
  NOR2_X1 U326 ( .A1(n124), .A2(n174), .ZN(ab_5__8_) );
  NOR2_X1 U327 ( .A1(n126), .A2(n174), .ZN(ab_5__7_) );
  NOR2_X1 U328 ( .A1(n128), .A2(n174), .ZN(ab_5__6_) );
  NOR2_X1 U329 ( .A1(n130), .A2(n174), .ZN(ab_5__5_) );
  NOR2_X1 U330 ( .A1(n132), .A2(n174), .ZN(ab_5__4_) );
  NOR2_X1 U331 ( .A1(n134), .A2(n174), .ZN(ab_5__3_) );
  NOR2_X1 U332 ( .A1(n136), .A2(n174), .ZN(ab_5__2_) );
  NOR2_X1 U333 ( .A1(n94), .A2(n174), .ZN(ab_5__23_) );
  NOR2_X1 U334 ( .A1(n96), .A2(n174), .ZN(ab_5__22_) );
  NOR2_X1 U335 ( .A1(n98), .A2(n174), .ZN(ab_5__21_) );
  NOR2_X1 U336 ( .A1(n100), .A2(n174), .ZN(ab_5__20_) );
  NOR2_X1 U337 ( .A1(n203), .A2(n173), .ZN(ab_5__1_) );
  NOR2_X1 U338 ( .A1(n102), .A2(n173), .ZN(ab_5__19_) );
  NOR2_X1 U339 ( .A1(n104), .A2(n173), .ZN(ab_5__18_) );
  NOR2_X1 U340 ( .A1(n106), .A2(n173), .ZN(ab_5__17_) );
  NOR2_X1 U341 ( .A1(n108), .A2(n173), .ZN(ab_5__16_) );
  NOR2_X1 U342 ( .A1(n110), .A2(n173), .ZN(ab_5__15_) );
  NOR2_X1 U343 ( .A1(n112), .A2(n173), .ZN(ab_5__14_) );
  NOR2_X1 U344 ( .A1(n114), .A2(n173), .ZN(ab_5__13_) );
  NOR2_X1 U345 ( .A1(n116), .A2(n173), .ZN(ab_5__12_) );
  NOR2_X1 U346 ( .A1(n118), .A2(n173), .ZN(ab_5__11_) );
  NOR2_X1 U347 ( .A1(n120), .A2(n173), .ZN(ab_5__10_) );
  NOR2_X1 U348 ( .A1(n204), .A2(n173), .ZN(ab_5__0_) );
  NOR2_X1 U349 ( .A1(n122), .A2(n176), .ZN(ab_4__9_) );
  NOR2_X1 U350 ( .A1(n124), .A2(n176), .ZN(ab_4__8_) );
  NOR2_X1 U351 ( .A1(n126), .A2(n176), .ZN(ab_4__7_) );
  NOR2_X1 U352 ( .A1(n128), .A2(n176), .ZN(ab_4__6_) );
  NOR2_X1 U353 ( .A1(n130), .A2(n176), .ZN(ab_4__5_) );
  NOR2_X1 U354 ( .A1(n132), .A2(n176), .ZN(ab_4__4_) );
  NOR2_X1 U355 ( .A1(n134), .A2(n176), .ZN(ab_4__3_) );
  NOR2_X1 U356 ( .A1(n136), .A2(n176), .ZN(ab_4__2_) );
  NOR2_X1 U357 ( .A1(n94), .A2(n176), .ZN(ab_4__23_) );
  NOR2_X1 U358 ( .A1(n96), .A2(n176), .ZN(ab_4__22_) );
  NOR2_X1 U359 ( .A1(n98), .A2(n176), .ZN(ab_4__21_) );
  NOR2_X1 U360 ( .A1(n100), .A2(n176), .ZN(ab_4__20_) );
  NOR2_X1 U361 ( .A1(n203), .A2(n175), .ZN(ab_4__1_) );
  NOR2_X1 U362 ( .A1(n102), .A2(n175), .ZN(ab_4__19_) );
  NOR2_X1 U363 ( .A1(n104), .A2(n175), .ZN(ab_4__18_) );
  NOR2_X1 U364 ( .A1(n106), .A2(n175), .ZN(ab_4__17_) );
  NOR2_X1 U365 ( .A1(n108), .A2(n175), .ZN(ab_4__16_) );
  NOR2_X1 U366 ( .A1(n110), .A2(n175), .ZN(ab_4__15_) );
  NOR2_X1 U367 ( .A1(n112), .A2(n175), .ZN(ab_4__14_) );
  NOR2_X1 U368 ( .A1(n114), .A2(n175), .ZN(ab_4__13_) );
  NOR2_X1 U369 ( .A1(n116), .A2(n175), .ZN(ab_4__12_) );
  NOR2_X1 U370 ( .A1(n118), .A2(n175), .ZN(ab_4__11_) );
  NOR2_X1 U371 ( .A1(n120), .A2(n175), .ZN(ab_4__10_) );
  NOR2_X1 U372 ( .A1(n204), .A2(n175), .ZN(ab_4__0_) );
  NOR2_X1 U373 ( .A1(n122), .A2(n178), .ZN(ab_3__9_) );
  NOR2_X1 U374 ( .A1(n124), .A2(n178), .ZN(ab_3__8_) );
  NOR2_X1 U375 ( .A1(n126), .A2(n178), .ZN(ab_3__7_) );
  NOR2_X1 U376 ( .A1(n128), .A2(n178), .ZN(ab_3__6_) );
  NOR2_X1 U377 ( .A1(n130), .A2(n178), .ZN(ab_3__5_) );
  NOR2_X1 U378 ( .A1(n132), .A2(n178), .ZN(ab_3__4_) );
  NOR2_X1 U379 ( .A1(n134), .A2(n178), .ZN(ab_3__3_) );
  NOR2_X1 U380 ( .A1(n136), .A2(n178), .ZN(ab_3__2_) );
  NOR2_X1 U381 ( .A1(n94), .A2(n178), .ZN(ab_3__23_) );
  NOR2_X1 U382 ( .A1(n96), .A2(n178), .ZN(ab_3__22_) );
  NOR2_X1 U383 ( .A1(n98), .A2(n178), .ZN(ab_3__21_) );
  NOR2_X1 U384 ( .A1(n100), .A2(n178), .ZN(ab_3__20_) );
  NOR2_X1 U385 ( .A1(n203), .A2(n177), .ZN(ab_3__1_) );
  NOR2_X1 U386 ( .A1(n102), .A2(n177), .ZN(ab_3__19_) );
  NOR2_X1 U387 ( .A1(n104), .A2(n177), .ZN(ab_3__18_) );
  NOR2_X1 U388 ( .A1(n106), .A2(n177), .ZN(ab_3__17_) );
  NOR2_X1 U389 ( .A1(n108), .A2(n177), .ZN(ab_3__16_) );
  NOR2_X1 U390 ( .A1(n110), .A2(n177), .ZN(ab_3__15_) );
  NOR2_X1 U391 ( .A1(n112), .A2(n177), .ZN(ab_3__14_) );
  NOR2_X1 U392 ( .A1(n114), .A2(n177), .ZN(ab_3__13_) );
  NOR2_X1 U393 ( .A1(n116), .A2(n177), .ZN(ab_3__12_) );
  NOR2_X1 U394 ( .A1(n118), .A2(n177), .ZN(ab_3__11_) );
  NOR2_X1 U395 ( .A1(n120), .A2(n177), .ZN(ab_3__10_) );
  NOR2_X1 U396 ( .A1(n204), .A2(n177), .ZN(ab_3__0_) );
  NOR2_X1 U397 ( .A1(n122), .A2(n180), .ZN(ab_2__9_) );
  NOR2_X1 U398 ( .A1(n124), .A2(n180), .ZN(ab_2__8_) );
  NOR2_X1 U399 ( .A1(n126), .A2(n180), .ZN(ab_2__7_) );
  NOR2_X1 U400 ( .A1(n128), .A2(n180), .ZN(ab_2__6_) );
  NOR2_X1 U401 ( .A1(n130), .A2(n180), .ZN(ab_2__5_) );
  NOR2_X1 U402 ( .A1(n132), .A2(n180), .ZN(ab_2__4_) );
  NOR2_X1 U403 ( .A1(n134), .A2(n180), .ZN(ab_2__3_) );
  NOR2_X1 U404 ( .A1(n136), .A2(n180), .ZN(ab_2__2_) );
  NOR2_X1 U405 ( .A1(n94), .A2(n180), .ZN(ab_2__23_) );
  NOR2_X1 U406 ( .A1(n96), .A2(n180), .ZN(ab_2__22_) );
  NOR2_X1 U407 ( .A1(n98), .A2(n180), .ZN(ab_2__21_) );
  NOR2_X1 U408 ( .A1(n100), .A2(n180), .ZN(ab_2__20_) );
  NOR2_X1 U409 ( .A1(n203), .A2(n179), .ZN(ab_2__1_) );
  NOR2_X1 U410 ( .A1(n102), .A2(n179), .ZN(ab_2__19_) );
  NOR2_X1 U411 ( .A1(n104), .A2(n179), .ZN(ab_2__18_) );
  NOR2_X1 U412 ( .A1(n106), .A2(n179), .ZN(ab_2__17_) );
  NOR2_X1 U413 ( .A1(n108), .A2(n179), .ZN(ab_2__16_) );
  NOR2_X1 U414 ( .A1(n110), .A2(n179), .ZN(ab_2__15_) );
  NOR2_X1 U415 ( .A1(n112), .A2(n179), .ZN(ab_2__14_) );
  NOR2_X1 U416 ( .A1(n114), .A2(n179), .ZN(ab_2__13_) );
  NOR2_X1 U417 ( .A1(n116), .A2(n179), .ZN(ab_2__12_) );
  NOR2_X1 U418 ( .A1(n118), .A2(n179), .ZN(ab_2__11_) );
  NOR2_X1 U419 ( .A1(n120), .A2(n179), .ZN(ab_2__10_) );
  NOR2_X1 U420 ( .A1(n204), .A2(n179), .ZN(ab_2__0_) );
  NOR2_X1 U421 ( .A1(n122), .A2(n138), .ZN(ab_23__9_) );
  NOR2_X1 U422 ( .A1(n124), .A2(n138), .ZN(ab_23__8_) );
  NOR2_X1 U423 ( .A1(n126), .A2(n138), .ZN(ab_23__7_) );
  NOR2_X1 U424 ( .A1(n128), .A2(n138), .ZN(ab_23__6_) );
  NOR2_X1 U425 ( .A1(n130), .A2(n138), .ZN(ab_23__5_) );
  NOR2_X1 U426 ( .A1(n132), .A2(n138), .ZN(ab_23__4_) );
  NOR2_X1 U427 ( .A1(n134), .A2(n138), .ZN(ab_23__3_) );
  NOR2_X1 U428 ( .A1(n136), .A2(n138), .ZN(ab_23__2_) );
  NOR2_X1 U429 ( .A1(n94), .A2(n138), .ZN(ab_23__23_) );
  NOR2_X1 U430 ( .A1(n96), .A2(n138), .ZN(ab_23__22_) );
  NOR2_X1 U431 ( .A1(n98), .A2(n138), .ZN(ab_23__21_) );
  NOR2_X1 U432 ( .A1(n100), .A2(n138), .ZN(ab_23__20_) );
  NOR2_X1 U433 ( .A1(n203), .A2(n137), .ZN(ab_23__1_) );
  NOR2_X1 U434 ( .A1(n102), .A2(n137), .ZN(ab_23__19_) );
  NOR2_X1 U435 ( .A1(n104), .A2(n137), .ZN(ab_23__18_) );
  NOR2_X1 U436 ( .A1(n106), .A2(n137), .ZN(ab_23__17_) );
  NOR2_X1 U437 ( .A1(n108), .A2(n137), .ZN(ab_23__16_) );
  NOR2_X1 U438 ( .A1(n110), .A2(n137), .ZN(ab_23__15_) );
  NOR2_X1 U439 ( .A1(n112), .A2(n137), .ZN(ab_23__14_) );
  NOR2_X1 U440 ( .A1(n114), .A2(n137), .ZN(ab_23__13_) );
  NOR2_X1 U441 ( .A1(n116), .A2(n137), .ZN(ab_23__12_) );
  NOR2_X1 U442 ( .A1(n118), .A2(n137), .ZN(ab_23__11_) );
  NOR2_X1 U443 ( .A1(n120), .A2(n137), .ZN(ab_23__10_) );
  NOR2_X1 U444 ( .A1(n204), .A2(n137), .ZN(ab_23__0_) );
  NOR2_X1 U445 ( .A1(n122), .A2(n140), .ZN(ab_22__9_) );
  NOR2_X1 U446 ( .A1(n124), .A2(n140), .ZN(ab_22__8_) );
  NOR2_X1 U447 ( .A1(n126), .A2(n140), .ZN(ab_22__7_) );
  NOR2_X1 U448 ( .A1(n128), .A2(n140), .ZN(ab_22__6_) );
  NOR2_X1 U449 ( .A1(n130), .A2(n140), .ZN(ab_22__5_) );
  NOR2_X1 U450 ( .A1(n132), .A2(n140), .ZN(ab_22__4_) );
  NOR2_X1 U451 ( .A1(n134), .A2(n140), .ZN(ab_22__3_) );
  NOR2_X1 U452 ( .A1(n136), .A2(n140), .ZN(ab_22__2_) );
  NOR2_X1 U453 ( .A1(n94), .A2(n140), .ZN(ab_22__23_) );
  NOR2_X1 U454 ( .A1(n96), .A2(n140), .ZN(ab_22__22_) );
  NOR2_X1 U455 ( .A1(n98), .A2(n140), .ZN(ab_22__21_) );
  NOR2_X1 U456 ( .A1(n100), .A2(n140), .ZN(ab_22__20_) );
  NOR2_X1 U457 ( .A1(n203), .A2(n139), .ZN(ab_22__1_) );
  NOR2_X1 U458 ( .A1(n102), .A2(n139), .ZN(ab_22__19_) );
  NOR2_X1 U459 ( .A1(n104), .A2(n139), .ZN(ab_22__18_) );
  NOR2_X1 U460 ( .A1(n106), .A2(n139), .ZN(ab_22__17_) );
  NOR2_X1 U461 ( .A1(n108), .A2(n139), .ZN(ab_22__16_) );
  NOR2_X1 U462 ( .A1(n110), .A2(n139), .ZN(ab_22__15_) );
  NOR2_X1 U463 ( .A1(n112), .A2(n139), .ZN(ab_22__14_) );
  NOR2_X1 U464 ( .A1(n114), .A2(n139), .ZN(ab_22__13_) );
  NOR2_X1 U465 ( .A1(n116), .A2(n139), .ZN(ab_22__12_) );
  NOR2_X1 U466 ( .A1(n118), .A2(n139), .ZN(ab_22__11_) );
  NOR2_X1 U467 ( .A1(n120), .A2(n139), .ZN(ab_22__10_) );
  NOR2_X1 U468 ( .A1(n204), .A2(n139), .ZN(ab_22__0_) );
  NOR2_X1 U469 ( .A1(n122), .A2(n142), .ZN(ab_21__9_) );
  NOR2_X1 U470 ( .A1(n124), .A2(n142), .ZN(ab_21__8_) );
  NOR2_X1 U471 ( .A1(n126), .A2(n142), .ZN(ab_21__7_) );
  NOR2_X1 U472 ( .A1(n128), .A2(n142), .ZN(ab_21__6_) );
  NOR2_X1 U473 ( .A1(n130), .A2(n142), .ZN(ab_21__5_) );
  NOR2_X1 U474 ( .A1(n132), .A2(n142), .ZN(ab_21__4_) );
  NOR2_X1 U475 ( .A1(n134), .A2(n142), .ZN(ab_21__3_) );
  NOR2_X1 U476 ( .A1(n136), .A2(n142), .ZN(ab_21__2_) );
  NOR2_X1 U477 ( .A1(n94), .A2(n142), .ZN(ab_21__23_) );
  NOR2_X1 U478 ( .A1(n96), .A2(n142), .ZN(ab_21__22_) );
  NOR2_X1 U479 ( .A1(n98), .A2(n142), .ZN(ab_21__21_) );
  NOR2_X1 U480 ( .A1(n100), .A2(n142), .ZN(ab_21__20_) );
  NOR2_X1 U481 ( .A1(n203), .A2(n141), .ZN(ab_21__1_) );
  NOR2_X1 U482 ( .A1(n102), .A2(n141), .ZN(ab_21__19_) );
  NOR2_X1 U483 ( .A1(n104), .A2(n141), .ZN(ab_21__18_) );
  NOR2_X1 U484 ( .A1(n106), .A2(n141), .ZN(ab_21__17_) );
  NOR2_X1 U485 ( .A1(n108), .A2(n141), .ZN(ab_21__16_) );
  NOR2_X1 U486 ( .A1(n110), .A2(n141), .ZN(ab_21__15_) );
  NOR2_X1 U487 ( .A1(n112), .A2(n141), .ZN(ab_21__14_) );
  NOR2_X1 U488 ( .A1(n114), .A2(n141), .ZN(ab_21__13_) );
  NOR2_X1 U489 ( .A1(n116), .A2(n141), .ZN(ab_21__12_) );
  NOR2_X1 U490 ( .A1(n118), .A2(n141), .ZN(ab_21__11_) );
  NOR2_X1 U491 ( .A1(n120), .A2(n141), .ZN(ab_21__10_) );
  NOR2_X1 U492 ( .A1(n204), .A2(n141), .ZN(ab_21__0_) );
  NOR2_X1 U493 ( .A1(n122), .A2(n144), .ZN(ab_20__9_) );
  NOR2_X1 U494 ( .A1(n124), .A2(n144), .ZN(ab_20__8_) );
  NOR2_X1 U495 ( .A1(n126), .A2(n144), .ZN(ab_20__7_) );
  NOR2_X1 U496 ( .A1(n128), .A2(n144), .ZN(ab_20__6_) );
  NOR2_X1 U497 ( .A1(n130), .A2(n144), .ZN(ab_20__5_) );
  NOR2_X1 U498 ( .A1(n132), .A2(n144), .ZN(ab_20__4_) );
  NOR2_X1 U499 ( .A1(n134), .A2(n144), .ZN(ab_20__3_) );
  NOR2_X1 U500 ( .A1(n136), .A2(n144), .ZN(ab_20__2_) );
  NOR2_X1 U501 ( .A1(n94), .A2(n144), .ZN(ab_20__23_) );
  NOR2_X1 U502 ( .A1(n96), .A2(n144), .ZN(ab_20__22_) );
  NOR2_X1 U503 ( .A1(n98), .A2(n144), .ZN(ab_20__21_) );
  NOR2_X1 U504 ( .A1(n100), .A2(n144), .ZN(ab_20__20_) );
  NOR2_X1 U505 ( .A1(n203), .A2(n143), .ZN(ab_20__1_) );
  NOR2_X1 U506 ( .A1(n102), .A2(n143), .ZN(ab_20__19_) );
  NOR2_X1 U507 ( .A1(n104), .A2(n143), .ZN(ab_20__18_) );
  NOR2_X1 U508 ( .A1(n106), .A2(n143), .ZN(ab_20__17_) );
  NOR2_X1 U509 ( .A1(n108), .A2(n143), .ZN(ab_20__16_) );
  NOR2_X1 U510 ( .A1(n110), .A2(n143), .ZN(ab_20__15_) );
  NOR2_X1 U511 ( .A1(n112), .A2(n143), .ZN(ab_20__14_) );
  NOR2_X1 U512 ( .A1(n114), .A2(n143), .ZN(ab_20__13_) );
  NOR2_X1 U513 ( .A1(n116), .A2(n143), .ZN(ab_20__12_) );
  NOR2_X1 U514 ( .A1(n118), .A2(n143), .ZN(ab_20__11_) );
  NOR2_X1 U515 ( .A1(n120), .A2(n143), .ZN(ab_20__10_) );
  NOR2_X1 U516 ( .A1(n204), .A2(n143), .ZN(ab_20__0_) );
  NOR2_X1 U517 ( .A1(n121), .A2(n227), .ZN(ab_1__9_) );
  NOR2_X1 U518 ( .A1(n123), .A2(n227), .ZN(ab_1__8_) );
  NOR2_X1 U519 ( .A1(n125), .A2(n227), .ZN(ab_1__7_) );
  NOR2_X1 U520 ( .A1(n127), .A2(n227), .ZN(ab_1__6_) );
  NOR2_X1 U521 ( .A1(n129), .A2(n227), .ZN(ab_1__5_) );
  NOR2_X1 U522 ( .A1(n131), .A2(n227), .ZN(ab_1__4_) );
  NOR2_X1 U523 ( .A1(n133), .A2(n227), .ZN(ab_1__3_) );
  NOR2_X1 U524 ( .A1(n135), .A2(n227), .ZN(ab_1__2_) );
  NOR2_X1 U525 ( .A1(n93), .A2(n227), .ZN(ab_1__23_) );
  NOR2_X1 U526 ( .A1(n95), .A2(n227), .ZN(ab_1__22_) );
  NOR2_X1 U527 ( .A1(n97), .A2(n227), .ZN(ab_1__21_) );
  NOR2_X1 U528 ( .A1(n99), .A2(n227), .ZN(ab_1__20_) );
  NOR2_X1 U529 ( .A1(n101), .A2(n227), .ZN(ab_1__19_) );
  NOR2_X1 U530 ( .A1(n103), .A2(n227), .ZN(ab_1__18_) );
  NOR2_X1 U531 ( .A1(n105), .A2(n227), .ZN(ab_1__17_) );
  NOR2_X1 U532 ( .A1(n107), .A2(n227), .ZN(ab_1__16_) );
  NOR2_X1 U533 ( .A1(n109), .A2(n227), .ZN(ab_1__15_) );
  NOR2_X1 U534 ( .A1(n111), .A2(n227), .ZN(ab_1__14_) );
  NOR2_X1 U535 ( .A1(n113), .A2(n227), .ZN(ab_1__13_) );
  NOR2_X1 U536 ( .A1(n115), .A2(n227), .ZN(ab_1__12_) );
  NOR2_X1 U537 ( .A1(n117), .A2(n227), .ZN(ab_1__11_) );
  NOR2_X1 U538 ( .A1(n119), .A2(n227), .ZN(ab_1__10_) );
  NOR2_X1 U539 ( .A1(n121), .A2(n146), .ZN(ab_19__9_) );
  NOR2_X1 U540 ( .A1(n123), .A2(n146), .ZN(ab_19__8_) );
  NOR2_X1 U541 ( .A1(n125), .A2(n146), .ZN(ab_19__7_) );
  NOR2_X1 U542 ( .A1(n127), .A2(n146), .ZN(ab_19__6_) );
  NOR2_X1 U543 ( .A1(n129), .A2(n146), .ZN(ab_19__5_) );
  NOR2_X1 U544 ( .A1(n131), .A2(n146), .ZN(ab_19__4_) );
  NOR2_X1 U545 ( .A1(n133), .A2(n146), .ZN(ab_19__3_) );
  NOR2_X1 U546 ( .A1(n135), .A2(n146), .ZN(ab_19__2_) );
  NOR2_X1 U547 ( .A1(n93), .A2(n146), .ZN(ab_19__23_) );
  NOR2_X1 U548 ( .A1(n95), .A2(n146), .ZN(ab_19__22_) );
  NOR2_X1 U549 ( .A1(n97), .A2(n146), .ZN(ab_19__21_) );
  NOR2_X1 U550 ( .A1(n99), .A2(n146), .ZN(ab_19__20_) );
  NOR2_X1 U551 ( .A1(n203), .A2(n145), .ZN(ab_19__1_) );
  NOR2_X1 U552 ( .A1(n101), .A2(n145), .ZN(ab_19__19_) );
  NOR2_X1 U553 ( .A1(n103), .A2(n145), .ZN(ab_19__18_) );
  NOR2_X1 U554 ( .A1(n105), .A2(n145), .ZN(ab_19__17_) );
  NOR2_X1 U555 ( .A1(n107), .A2(n145), .ZN(ab_19__16_) );
  NOR2_X1 U556 ( .A1(n109), .A2(n145), .ZN(ab_19__15_) );
  NOR2_X1 U557 ( .A1(n111), .A2(n145), .ZN(ab_19__14_) );
  NOR2_X1 U558 ( .A1(n113), .A2(n145), .ZN(ab_19__13_) );
  NOR2_X1 U559 ( .A1(n115), .A2(n145), .ZN(ab_19__12_) );
  NOR2_X1 U560 ( .A1(n117), .A2(n145), .ZN(ab_19__11_) );
  NOR2_X1 U561 ( .A1(n119), .A2(n145), .ZN(ab_19__10_) );
  NOR2_X1 U562 ( .A1(n204), .A2(n145), .ZN(ab_19__0_) );
  NOR2_X1 U563 ( .A1(n121), .A2(n148), .ZN(ab_18__9_) );
  NOR2_X1 U564 ( .A1(n123), .A2(n148), .ZN(ab_18__8_) );
  NOR2_X1 U565 ( .A1(n125), .A2(n148), .ZN(ab_18__7_) );
  NOR2_X1 U566 ( .A1(n127), .A2(n148), .ZN(ab_18__6_) );
  NOR2_X1 U567 ( .A1(n129), .A2(n148), .ZN(ab_18__5_) );
  NOR2_X1 U568 ( .A1(n131), .A2(n148), .ZN(ab_18__4_) );
  NOR2_X1 U569 ( .A1(n133), .A2(n148), .ZN(ab_18__3_) );
  NOR2_X1 U570 ( .A1(n135), .A2(n148), .ZN(ab_18__2_) );
  NOR2_X1 U571 ( .A1(n93), .A2(n148), .ZN(ab_18__23_) );
  NOR2_X1 U572 ( .A1(n95), .A2(n148), .ZN(ab_18__22_) );
  NOR2_X1 U573 ( .A1(n97), .A2(n148), .ZN(ab_18__21_) );
  NOR2_X1 U574 ( .A1(n99), .A2(n148), .ZN(ab_18__20_) );
  NOR2_X1 U575 ( .A1(n203), .A2(n147), .ZN(ab_18__1_) );
  NOR2_X1 U576 ( .A1(n101), .A2(n147), .ZN(ab_18__19_) );
  NOR2_X1 U577 ( .A1(n103), .A2(n147), .ZN(ab_18__18_) );
  NOR2_X1 U578 ( .A1(n105), .A2(n147), .ZN(ab_18__17_) );
  NOR2_X1 U579 ( .A1(n107), .A2(n147), .ZN(ab_18__16_) );
  NOR2_X1 U580 ( .A1(n109), .A2(n147), .ZN(ab_18__15_) );
  NOR2_X1 U581 ( .A1(n111), .A2(n147), .ZN(ab_18__14_) );
  NOR2_X1 U582 ( .A1(n113), .A2(n147), .ZN(ab_18__13_) );
  NOR2_X1 U583 ( .A1(n115), .A2(n147), .ZN(ab_18__12_) );
  NOR2_X1 U584 ( .A1(n117), .A2(n147), .ZN(ab_18__11_) );
  NOR2_X1 U585 ( .A1(n119), .A2(n147), .ZN(ab_18__10_) );
  NOR2_X1 U586 ( .A1(n204), .A2(n147), .ZN(ab_18__0_) );
  NOR2_X1 U587 ( .A1(n121), .A2(n150), .ZN(ab_17__9_) );
  NOR2_X1 U588 ( .A1(n123), .A2(n150), .ZN(ab_17__8_) );
  NOR2_X1 U589 ( .A1(n125), .A2(n150), .ZN(ab_17__7_) );
  NOR2_X1 U590 ( .A1(n127), .A2(n150), .ZN(ab_17__6_) );
  NOR2_X1 U591 ( .A1(n129), .A2(n150), .ZN(ab_17__5_) );
  NOR2_X1 U592 ( .A1(n131), .A2(n150), .ZN(ab_17__4_) );
  NOR2_X1 U593 ( .A1(n133), .A2(n150), .ZN(ab_17__3_) );
  NOR2_X1 U594 ( .A1(n135), .A2(n150), .ZN(ab_17__2_) );
  NOR2_X1 U595 ( .A1(n93), .A2(n150), .ZN(ab_17__23_) );
  NOR2_X1 U596 ( .A1(n95), .A2(n150), .ZN(ab_17__22_) );
  NOR2_X1 U597 ( .A1(n97), .A2(n150), .ZN(ab_17__21_) );
  NOR2_X1 U598 ( .A1(n99), .A2(n150), .ZN(ab_17__20_) );
  NOR2_X1 U599 ( .A1(n203), .A2(n149), .ZN(ab_17__1_) );
  NOR2_X1 U600 ( .A1(n101), .A2(n149), .ZN(ab_17__19_) );
  NOR2_X1 U601 ( .A1(n103), .A2(n149), .ZN(ab_17__18_) );
  NOR2_X1 U602 ( .A1(n105), .A2(n149), .ZN(ab_17__17_) );
  NOR2_X1 U603 ( .A1(n107), .A2(n149), .ZN(ab_17__16_) );
  NOR2_X1 U604 ( .A1(n109), .A2(n149), .ZN(ab_17__15_) );
  NOR2_X1 U605 ( .A1(n111), .A2(n149), .ZN(ab_17__14_) );
  NOR2_X1 U606 ( .A1(n113), .A2(n149), .ZN(ab_17__13_) );
  NOR2_X1 U607 ( .A1(n115), .A2(n149), .ZN(ab_17__12_) );
  NOR2_X1 U608 ( .A1(n117), .A2(n149), .ZN(ab_17__11_) );
  NOR2_X1 U609 ( .A1(n119), .A2(n149), .ZN(ab_17__10_) );
  NOR2_X1 U610 ( .A1(n204), .A2(n149), .ZN(ab_17__0_) );
  NOR2_X1 U611 ( .A1(n121), .A2(n152), .ZN(ab_16__9_) );
  NOR2_X1 U612 ( .A1(n123), .A2(n152), .ZN(ab_16__8_) );
  NOR2_X1 U613 ( .A1(n125), .A2(n152), .ZN(ab_16__7_) );
  NOR2_X1 U614 ( .A1(n127), .A2(n152), .ZN(ab_16__6_) );
  NOR2_X1 U615 ( .A1(n129), .A2(n152), .ZN(ab_16__5_) );
  NOR2_X1 U616 ( .A1(n131), .A2(n152), .ZN(ab_16__4_) );
  NOR2_X1 U617 ( .A1(n133), .A2(n152), .ZN(ab_16__3_) );
  NOR2_X1 U618 ( .A1(n135), .A2(n152), .ZN(ab_16__2_) );
  NOR2_X1 U619 ( .A1(n93), .A2(n152), .ZN(ab_16__23_) );
  NOR2_X1 U620 ( .A1(n95), .A2(n152), .ZN(ab_16__22_) );
  NOR2_X1 U621 ( .A1(n97), .A2(n152), .ZN(ab_16__21_) );
  NOR2_X1 U622 ( .A1(n99), .A2(n152), .ZN(ab_16__20_) );
  NOR2_X1 U623 ( .A1(n203), .A2(n151), .ZN(ab_16__1_) );
  NOR2_X1 U624 ( .A1(n101), .A2(n151), .ZN(ab_16__19_) );
  NOR2_X1 U625 ( .A1(n103), .A2(n151), .ZN(ab_16__18_) );
  NOR2_X1 U626 ( .A1(n105), .A2(n151), .ZN(ab_16__17_) );
  NOR2_X1 U627 ( .A1(n107), .A2(n151), .ZN(ab_16__16_) );
  NOR2_X1 U628 ( .A1(n109), .A2(n151), .ZN(ab_16__15_) );
  NOR2_X1 U629 ( .A1(n111), .A2(n151), .ZN(ab_16__14_) );
  NOR2_X1 U630 ( .A1(n113), .A2(n151), .ZN(ab_16__13_) );
  NOR2_X1 U631 ( .A1(n115), .A2(n151), .ZN(ab_16__12_) );
  NOR2_X1 U632 ( .A1(n117), .A2(n151), .ZN(ab_16__11_) );
  NOR2_X1 U633 ( .A1(n119), .A2(n151), .ZN(ab_16__10_) );
  NOR2_X1 U634 ( .A1(n204), .A2(n151), .ZN(ab_16__0_) );
  NOR2_X1 U635 ( .A1(n121), .A2(n154), .ZN(ab_15__9_) );
  NOR2_X1 U636 ( .A1(n123), .A2(n154), .ZN(ab_15__8_) );
  NOR2_X1 U637 ( .A1(n125), .A2(n154), .ZN(ab_15__7_) );
  NOR2_X1 U638 ( .A1(n127), .A2(n154), .ZN(ab_15__6_) );
  NOR2_X1 U639 ( .A1(n129), .A2(n154), .ZN(ab_15__5_) );
  NOR2_X1 U640 ( .A1(n131), .A2(n154), .ZN(ab_15__4_) );
  NOR2_X1 U641 ( .A1(n133), .A2(n154), .ZN(ab_15__3_) );
  NOR2_X1 U642 ( .A1(n135), .A2(n154), .ZN(ab_15__2_) );
  NOR2_X1 U643 ( .A1(n93), .A2(n154), .ZN(ab_15__23_) );
  NOR2_X1 U644 ( .A1(n95), .A2(n154), .ZN(ab_15__22_) );
  NOR2_X1 U645 ( .A1(n97), .A2(n154), .ZN(ab_15__21_) );
  NOR2_X1 U646 ( .A1(n99), .A2(n154), .ZN(ab_15__20_) );
  NOR2_X1 U647 ( .A1(n203), .A2(n153), .ZN(ab_15__1_) );
  NOR2_X1 U648 ( .A1(n101), .A2(n153), .ZN(ab_15__19_) );
  NOR2_X1 U649 ( .A1(n103), .A2(n153), .ZN(ab_15__18_) );
  NOR2_X1 U650 ( .A1(n105), .A2(n153), .ZN(ab_15__17_) );
  NOR2_X1 U651 ( .A1(n107), .A2(n153), .ZN(ab_15__16_) );
  NOR2_X1 U652 ( .A1(n109), .A2(n153), .ZN(ab_15__15_) );
  NOR2_X1 U653 ( .A1(n111), .A2(n153), .ZN(ab_15__14_) );
  NOR2_X1 U654 ( .A1(n113), .A2(n153), .ZN(ab_15__13_) );
  NOR2_X1 U655 ( .A1(n115), .A2(n153), .ZN(ab_15__12_) );
  NOR2_X1 U656 ( .A1(n117), .A2(n153), .ZN(ab_15__11_) );
  NOR2_X1 U657 ( .A1(n119), .A2(n153), .ZN(ab_15__10_) );
  NOR2_X1 U658 ( .A1(n204), .A2(n153), .ZN(ab_15__0_) );
  NOR2_X1 U659 ( .A1(n121), .A2(n156), .ZN(ab_14__9_) );
  NOR2_X1 U660 ( .A1(n123), .A2(n156), .ZN(ab_14__8_) );
  NOR2_X1 U661 ( .A1(n125), .A2(n156), .ZN(ab_14__7_) );
  NOR2_X1 U662 ( .A1(n127), .A2(n156), .ZN(ab_14__6_) );
  NOR2_X1 U663 ( .A1(n129), .A2(n156), .ZN(ab_14__5_) );
  NOR2_X1 U664 ( .A1(n131), .A2(n156), .ZN(ab_14__4_) );
  NOR2_X1 U665 ( .A1(n133), .A2(n156), .ZN(ab_14__3_) );
  NOR2_X1 U666 ( .A1(n135), .A2(n156), .ZN(ab_14__2_) );
  NOR2_X1 U667 ( .A1(n93), .A2(n156), .ZN(ab_14__23_) );
  NOR2_X1 U668 ( .A1(n95), .A2(n156), .ZN(ab_14__22_) );
  NOR2_X1 U669 ( .A1(n97), .A2(n156), .ZN(ab_14__21_) );
  NOR2_X1 U670 ( .A1(n99), .A2(n156), .ZN(ab_14__20_) );
  NOR2_X1 U671 ( .A1(n203), .A2(n155), .ZN(ab_14__1_) );
  NOR2_X1 U672 ( .A1(n101), .A2(n155), .ZN(ab_14__19_) );
  NOR2_X1 U673 ( .A1(n103), .A2(n155), .ZN(ab_14__18_) );
  NOR2_X1 U674 ( .A1(n105), .A2(n155), .ZN(ab_14__17_) );
  NOR2_X1 U675 ( .A1(n107), .A2(n155), .ZN(ab_14__16_) );
  NOR2_X1 U676 ( .A1(n109), .A2(n155), .ZN(ab_14__15_) );
  NOR2_X1 U677 ( .A1(n111), .A2(n155), .ZN(ab_14__14_) );
  NOR2_X1 U678 ( .A1(n113), .A2(n155), .ZN(ab_14__13_) );
  NOR2_X1 U679 ( .A1(n115), .A2(n155), .ZN(ab_14__12_) );
  NOR2_X1 U680 ( .A1(n117), .A2(n155), .ZN(ab_14__11_) );
  NOR2_X1 U681 ( .A1(n119), .A2(n155), .ZN(ab_14__10_) );
  NOR2_X1 U682 ( .A1(n204), .A2(n155), .ZN(ab_14__0_) );
  NOR2_X1 U683 ( .A1(n121), .A2(n158), .ZN(ab_13__9_) );
  NOR2_X1 U684 ( .A1(n123), .A2(n158), .ZN(ab_13__8_) );
  NOR2_X1 U685 ( .A1(n125), .A2(n158), .ZN(ab_13__7_) );
  NOR2_X1 U686 ( .A1(n127), .A2(n158), .ZN(ab_13__6_) );
  NOR2_X1 U687 ( .A1(n129), .A2(n158), .ZN(ab_13__5_) );
  NOR2_X1 U688 ( .A1(n131), .A2(n158), .ZN(ab_13__4_) );
  NOR2_X1 U689 ( .A1(n133), .A2(n158), .ZN(ab_13__3_) );
  NOR2_X1 U690 ( .A1(n135), .A2(n158), .ZN(ab_13__2_) );
  NOR2_X1 U691 ( .A1(n93), .A2(n158), .ZN(ab_13__23_) );
  NOR2_X1 U692 ( .A1(n95), .A2(n158), .ZN(ab_13__22_) );
  NOR2_X1 U693 ( .A1(n97), .A2(n158), .ZN(ab_13__21_) );
  NOR2_X1 U694 ( .A1(n99), .A2(n158), .ZN(ab_13__20_) );
  NOR2_X1 U695 ( .A1(n203), .A2(n157), .ZN(ab_13__1_) );
  NOR2_X1 U696 ( .A1(n101), .A2(n157), .ZN(ab_13__19_) );
  NOR2_X1 U697 ( .A1(n103), .A2(n157), .ZN(ab_13__18_) );
  NOR2_X1 U698 ( .A1(n105), .A2(n157), .ZN(ab_13__17_) );
  NOR2_X1 U699 ( .A1(n107), .A2(n157), .ZN(ab_13__16_) );
  NOR2_X1 U700 ( .A1(n109), .A2(n157), .ZN(ab_13__15_) );
  NOR2_X1 U701 ( .A1(n111), .A2(n157), .ZN(ab_13__14_) );
  NOR2_X1 U702 ( .A1(n113), .A2(n157), .ZN(ab_13__13_) );
  NOR2_X1 U703 ( .A1(n115), .A2(n157), .ZN(ab_13__12_) );
  NOR2_X1 U704 ( .A1(n117), .A2(n157), .ZN(ab_13__11_) );
  NOR2_X1 U705 ( .A1(n119), .A2(n157), .ZN(ab_13__10_) );
  NOR2_X1 U706 ( .A1(n204), .A2(n157), .ZN(ab_13__0_) );
  NOR2_X1 U707 ( .A1(n121), .A2(n160), .ZN(ab_12__9_) );
  NOR2_X1 U708 ( .A1(n123), .A2(n160), .ZN(ab_12__8_) );
  NOR2_X1 U709 ( .A1(n125), .A2(n160), .ZN(ab_12__7_) );
  NOR2_X1 U710 ( .A1(n127), .A2(n160), .ZN(ab_12__6_) );
  NOR2_X1 U711 ( .A1(n129), .A2(n160), .ZN(ab_12__5_) );
  NOR2_X1 U712 ( .A1(n131), .A2(n160), .ZN(ab_12__4_) );
  NOR2_X1 U713 ( .A1(n133), .A2(n160), .ZN(ab_12__3_) );
  NOR2_X1 U714 ( .A1(n135), .A2(n160), .ZN(ab_12__2_) );
  NOR2_X1 U715 ( .A1(n93), .A2(n160), .ZN(ab_12__23_) );
  NOR2_X1 U716 ( .A1(n95), .A2(n160), .ZN(ab_12__22_) );
  NOR2_X1 U717 ( .A1(n97), .A2(n160), .ZN(ab_12__21_) );
  NOR2_X1 U718 ( .A1(n99), .A2(n160), .ZN(ab_12__20_) );
  NOR2_X1 U719 ( .A1(n203), .A2(n159), .ZN(ab_12__1_) );
  NOR2_X1 U720 ( .A1(n101), .A2(n159), .ZN(ab_12__19_) );
  NOR2_X1 U721 ( .A1(n103), .A2(n159), .ZN(ab_12__18_) );
  NOR2_X1 U722 ( .A1(n105), .A2(n159), .ZN(ab_12__17_) );
  NOR2_X1 U723 ( .A1(n107), .A2(n159), .ZN(ab_12__16_) );
  NOR2_X1 U724 ( .A1(n109), .A2(n159), .ZN(ab_12__15_) );
  NOR2_X1 U725 ( .A1(n111), .A2(n159), .ZN(ab_12__14_) );
  NOR2_X1 U726 ( .A1(n113), .A2(n159), .ZN(ab_12__13_) );
  NOR2_X1 U727 ( .A1(n115), .A2(n159), .ZN(ab_12__12_) );
  NOR2_X1 U728 ( .A1(n117), .A2(n159), .ZN(ab_12__11_) );
  NOR2_X1 U729 ( .A1(n119), .A2(n159), .ZN(ab_12__10_) );
  NOR2_X1 U730 ( .A1(n204), .A2(n159), .ZN(ab_12__0_) );
  NOR2_X1 U731 ( .A1(n121), .A2(n162), .ZN(ab_11__9_) );
  NOR2_X1 U732 ( .A1(n123), .A2(n162), .ZN(ab_11__8_) );
  NOR2_X1 U733 ( .A1(n125), .A2(n162), .ZN(ab_11__7_) );
  NOR2_X1 U734 ( .A1(n127), .A2(n162), .ZN(ab_11__6_) );
  NOR2_X1 U735 ( .A1(n129), .A2(n162), .ZN(ab_11__5_) );
  NOR2_X1 U736 ( .A1(n131), .A2(n162), .ZN(ab_11__4_) );
  NOR2_X1 U737 ( .A1(n133), .A2(n162), .ZN(ab_11__3_) );
  NOR2_X1 U738 ( .A1(n135), .A2(n162), .ZN(ab_11__2_) );
  NOR2_X1 U739 ( .A1(n93), .A2(n162), .ZN(ab_11__23_) );
  NOR2_X1 U740 ( .A1(n95), .A2(n162), .ZN(ab_11__22_) );
  NOR2_X1 U741 ( .A1(n97), .A2(n162), .ZN(ab_11__21_) );
  NOR2_X1 U742 ( .A1(n99), .A2(n162), .ZN(ab_11__20_) );
  NOR2_X1 U743 ( .A1(n203), .A2(n161), .ZN(ab_11__1_) );
  NOR2_X1 U744 ( .A1(n101), .A2(n161), .ZN(ab_11__19_) );
  NOR2_X1 U745 ( .A1(n103), .A2(n161), .ZN(ab_11__18_) );
  NOR2_X1 U746 ( .A1(n105), .A2(n161), .ZN(ab_11__17_) );
  NOR2_X1 U747 ( .A1(n107), .A2(n161), .ZN(ab_11__16_) );
  NOR2_X1 U748 ( .A1(n109), .A2(n161), .ZN(ab_11__15_) );
  NOR2_X1 U749 ( .A1(n111), .A2(n161), .ZN(ab_11__14_) );
  NOR2_X1 U750 ( .A1(n113), .A2(n161), .ZN(ab_11__13_) );
  NOR2_X1 U751 ( .A1(n115), .A2(n161), .ZN(ab_11__12_) );
  NOR2_X1 U752 ( .A1(n117), .A2(n161), .ZN(ab_11__11_) );
  NOR2_X1 U753 ( .A1(n119), .A2(n161), .ZN(ab_11__10_) );
  NOR2_X1 U754 ( .A1(n204), .A2(n161), .ZN(ab_11__0_) );
  NOR2_X1 U755 ( .A1(n121), .A2(n164), .ZN(ab_10__9_) );
  NOR2_X1 U756 ( .A1(n123), .A2(n164), .ZN(ab_10__8_) );
  NOR2_X1 U757 ( .A1(n125), .A2(n164), .ZN(ab_10__7_) );
  NOR2_X1 U758 ( .A1(n127), .A2(n164), .ZN(ab_10__6_) );
  NOR2_X1 U759 ( .A1(n129), .A2(n164), .ZN(ab_10__5_) );
  NOR2_X1 U760 ( .A1(n131), .A2(n164), .ZN(ab_10__4_) );
  NOR2_X1 U761 ( .A1(n133), .A2(n164), .ZN(ab_10__3_) );
  NOR2_X1 U762 ( .A1(n135), .A2(n164), .ZN(ab_10__2_) );
  NOR2_X1 U763 ( .A1(n93), .A2(n164), .ZN(ab_10__23_) );
  NOR2_X1 U764 ( .A1(n95), .A2(n164), .ZN(ab_10__22_) );
  NOR2_X1 U765 ( .A1(n97), .A2(n164), .ZN(ab_10__21_) );
  NOR2_X1 U766 ( .A1(n99), .A2(n164), .ZN(ab_10__20_) );
  NOR2_X1 U767 ( .A1(n203), .A2(n163), .ZN(ab_10__1_) );
  NOR2_X1 U768 ( .A1(n101), .A2(n163), .ZN(ab_10__19_) );
  NOR2_X1 U769 ( .A1(n103), .A2(n163), .ZN(ab_10__18_) );
  NOR2_X1 U770 ( .A1(n105), .A2(n163), .ZN(ab_10__17_) );
  NOR2_X1 U771 ( .A1(n107), .A2(n163), .ZN(ab_10__16_) );
  NOR2_X1 U772 ( .A1(n109), .A2(n163), .ZN(ab_10__15_) );
  NOR2_X1 U773 ( .A1(n111), .A2(n163), .ZN(ab_10__14_) );
  NOR2_X1 U774 ( .A1(n113), .A2(n163), .ZN(ab_10__13_) );
  NOR2_X1 U775 ( .A1(n115), .A2(n163), .ZN(ab_10__12_) );
  NOR2_X1 U776 ( .A1(n117), .A2(n163), .ZN(ab_10__11_) );
  NOR2_X1 U777 ( .A1(n119), .A2(n163), .ZN(ab_10__10_) );
  NOR2_X1 U778 ( .A1(n204), .A2(n163), .ZN(ab_10__0_) );
  NOR2_X1 U779 ( .A1(n121), .A2(n228), .ZN(ab_0__9_) );
  NOR2_X1 U780 ( .A1(n123), .A2(n228), .ZN(ab_0__8_) );
  NOR2_X1 U781 ( .A1(n125), .A2(n228), .ZN(ab_0__7_) );
  NOR2_X1 U782 ( .A1(n127), .A2(n228), .ZN(ab_0__6_) );
  NOR2_X1 U783 ( .A1(n129), .A2(n228), .ZN(ab_0__5_) );
  NOR2_X1 U784 ( .A1(n131), .A2(n228), .ZN(ab_0__4_) );
  NOR2_X1 U785 ( .A1(n133), .A2(n228), .ZN(ab_0__3_) );
  NOR2_X1 U786 ( .A1(n135), .A2(n228), .ZN(ab_0__2_) );
  NOR2_X1 U787 ( .A1(n93), .A2(n228), .ZN(ab_0__23_) );
  NOR2_X1 U788 ( .A1(n95), .A2(n228), .ZN(ab_0__22_) );
  NOR2_X1 U789 ( .A1(n97), .A2(n228), .ZN(ab_0__21_) );
  NOR2_X1 U790 ( .A1(n99), .A2(n228), .ZN(ab_0__20_) );
  NOR2_X1 U791 ( .A1(n101), .A2(n228), .ZN(ab_0__19_) );
  NOR2_X1 U792 ( .A1(n103), .A2(n228), .ZN(ab_0__18_) );
  NOR2_X1 U793 ( .A1(n105), .A2(n228), .ZN(ab_0__17_) );
  NOR2_X1 U794 ( .A1(n107), .A2(n228), .ZN(ab_0__16_) );
  NOR2_X1 U795 ( .A1(n109), .A2(n228), .ZN(ab_0__15_) );
  NOR2_X1 U796 ( .A1(n111), .A2(n228), .ZN(ab_0__14_) );
  NOR2_X1 U797 ( .A1(n113), .A2(n228), .ZN(ab_0__13_) );
  NOR2_X1 U798 ( .A1(n115), .A2(n228), .ZN(ab_0__12_) );
  NOR2_X1 U799 ( .A1(n117), .A2(n228), .ZN(ab_0__11_) );
  NOR2_X1 U800 ( .A1(n119), .A2(n228), .ZN(ab_0__10_) );
  AND3_X1 U801 ( .A1(ab_1__1_), .A2(B[0]), .A3(A[0]), .ZN(CARRYB_1__0_) );
  NOR2_X1 U802 ( .A1(n227), .A2(n203), .ZN(ab_1__1_) );
endmodule


module fpMultiplier_DW01_add_1 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:2] carry;

  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(SUM[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(B[0]), .A2(A[0]), .ZN(n1) );
  XOR2_X1 U2 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module fpMultiplier ( clk, reset, enable, A, B, result, overflow );
  input [31:0] A;
  input [31:0] B;
  output [31:0] result;
  input clk, reset, enable;
  output overflow;
  wire   N27, n8, n9, n11, n141, n142, n143, n168, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, N90, N80,
         add_0_root_sub_1_root_add_24_2_carry_2_,
         add_0_root_sub_1_root_add_24_2_A_0_,
         add_0_root_sub_1_root_add_24_2_A_1_,
         add_0_root_sub_1_root_add_24_2_A_2_,
         add_0_root_sub_1_root_add_24_2_A_3_,
         add_0_root_sub_1_root_add_24_2_A_4_,
         add_0_root_sub_1_root_add_24_2_A_5_,
         add_0_root_sub_1_root_add_24_2_A_6_,
         add_0_root_sub_1_root_add_24_2_A_7_,
         add_0_root_sub_1_root_add_24_2_A_8_, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, SYNOPSYS_UNCONNECTED_1,
         SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3,
         SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5,
         SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7,
         SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9,
         SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11,
         SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13,
         SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15,
         SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17,
         SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19,
         SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21,
         SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23;
  wire   [30:23] regA;
  wire   [30:23] regB;
  wire   [23:0] MA;
  wire   [23:0] MB;
  wire   [46:23] mantissasProduct;

  DFF_X1 result_reg_31_ ( .D(n267), .CK(clk), .Q(result[31]), .QN(n202) );
  DFF_X1 result_reg_30_ ( .D(n266), .CK(clk), .Q(result[30]), .QN(n203) );
  DFF_X1 result_reg_29_ ( .D(n265), .CK(clk), .Q(result[29]), .QN(n204) );
  DFF_X1 result_reg_28_ ( .D(n264), .CK(clk), .Q(result[28]), .QN(n205) );
  DFF_X1 result_reg_27_ ( .D(n263), .CK(clk), .Q(result[27]), .QN(n206) );
  DFF_X1 result_reg_26_ ( .D(n262), .CK(clk), .Q(result[26]), .QN(n207) );
  DFF_X1 result_reg_25_ ( .D(n261), .CK(clk), .Q(result[25]), .QN(n208) );
  DFF_X1 result_reg_24_ ( .D(n260), .CK(clk), .Q(result[24]), .QN(n209) );
  DFF_X1 result_reg_23_ ( .D(n259), .CK(clk), .Q(result[23]), .QN(n210) );
  DFF_X1 result_reg_22_ ( .D(n258), .CK(clk), .Q(result[22]), .QN(n211) );
  DFF_X1 result_reg_21_ ( .D(n257), .CK(clk), .Q(result[21]), .QN(n212) );
  DFF_X1 result_reg_20_ ( .D(n256), .CK(clk), .Q(result[20]), .QN(n213) );
  DFF_X1 result_reg_19_ ( .D(n255), .CK(clk), .Q(result[19]), .QN(n214) );
  DFF_X1 result_reg_18_ ( .D(n254), .CK(clk), .Q(result[18]), .QN(n215) );
  DFF_X1 result_reg_17_ ( .D(n253), .CK(clk), .Q(result[17]), .QN(n216) );
  DFF_X1 result_reg_16_ ( .D(n252), .CK(clk), .Q(result[16]), .QN(n217) );
  DFF_X1 result_reg_15_ ( .D(n251), .CK(clk), .Q(result[15]), .QN(n218) );
  DFF_X1 result_reg_14_ ( .D(n250), .CK(clk), .Q(result[14]), .QN(n219) );
  DFF_X1 result_reg_13_ ( .D(n249), .CK(clk), .Q(result[13]), .QN(n220) );
  DFF_X1 result_reg_12_ ( .D(n248), .CK(clk), .Q(result[12]), .QN(n221) );
  DFF_X1 result_reg_11_ ( .D(n247), .CK(clk), .Q(result[11]), .QN(n222) );
  DFF_X1 result_reg_10_ ( .D(n246), .CK(clk), .Q(result[10]), .QN(n223) );
  DFF_X1 result_reg_9_ ( .D(n245), .CK(clk), .Q(result[9]), .QN(n224) );
  DFF_X1 result_reg_8_ ( .D(n244), .CK(clk), .Q(result[8]), .QN(n225) );
  DFF_X1 result_reg_7_ ( .D(n243), .CK(clk), .Q(result[7]), .QN(n226) );
  DFF_X1 result_reg_6_ ( .D(n242), .CK(clk), .Q(result[6]), .QN(n227) );
  DFF_X1 result_reg_5_ ( .D(n241), .CK(clk), .Q(result[5]), .QN(n228) );
  DFF_X1 result_reg_4_ ( .D(n240), .CK(clk), .Q(result[4]), .QN(n229) );
  DFF_X1 result_reg_3_ ( .D(n239), .CK(clk), .Q(result[3]), .QN(n230) );
  DFF_X1 result_reg_2_ ( .D(n238), .CK(clk), .Q(result[2]), .QN(n231) );
  DFF_X1 result_reg_1_ ( .D(n237), .CK(clk), .Q(result[1]), .QN(n232) );
  DFF_X1 result_reg_0_ ( .D(n236), .CK(clk), .Q(result[0]), .QN(n233) );
  DFF_X1 overflow_reg ( .D(n235), .CK(clk), .Q(overflow), .QN(n234) );
  fpMultiplier_DW02_mult_0 mult_21 ( .A(MA), .B(MB), .TC(1'b0), .PRODUCT({N90, 
        mantissasProduct, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, 
        SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, 
        SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, 
        SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10, 
        SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12, 
        SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14, 
        SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16, 
        SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18, 
        SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20, 
        SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22, 
        SYNOPSYS_UNCONNECTED_23}) );
  fpMultiplier_DW01_add_1 add_2_root_sub_1_root_add_24_2 ( .A({1'b0, regB}), 
        .B({1'b0, regA}), .CI(1'b0), .SUM({add_0_root_sub_1_root_add_24_2_A_8_, 
        add_0_root_sub_1_root_add_24_2_A_7_, 
        add_0_root_sub_1_root_add_24_2_A_6_, 
        add_0_root_sub_1_root_add_24_2_A_5_, 
        add_0_root_sub_1_root_add_24_2_A_4_, 
        add_0_root_sub_1_root_add_24_2_A_3_, 
        add_0_root_sub_1_root_add_24_2_A_2_, 
        add_0_root_sub_1_root_add_24_2_A_1_, 
        add_0_root_sub_1_root_add_24_2_A_0_}) );
  FA_X1 add_0_root_sub_1_root_add_24_2_U1_1 ( .A(
        add_0_root_sub_1_root_add_24_2_A_1_), .B(N90), .CI(n340), .CO(
        add_0_root_sub_1_root_add_24_2_carry_2_), .S(N27) );
  DFF_X1 regB_reg_31_ ( .D(n331), .CK(clk), .Q(n201), .QN(n455) );
  DFF_X1 regB_reg_30_ ( .D(n330), .CK(clk), .Q(regB[30]), .QN(n456) );
  DFF_X1 regB_reg_29_ ( .D(n329), .CK(clk), .Q(regB[29]), .QN(n457) );
  DFF_X1 regB_reg_28_ ( .D(n328), .CK(clk), .Q(regB[28]), .QN(n458) );
  DFF_X1 regB_reg_27_ ( .D(n327), .CK(clk), .Q(regB[27]), .QN(n459) );
  DFF_X1 regB_reg_26_ ( .D(n326), .CK(clk), .Q(regB[26]), .QN(n460) );
  DFF_X1 regB_reg_25_ ( .D(n325), .CK(clk), .Q(regB[25]), .QN(n461) );
  DFF_X1 regB_reg_24_ ( .D(n324), .CK(clk), .Q(regB[24]), .QN(n462) );
  DFF_X1 regB_reg_23_ ( .D(n323), .CK(clk), .Q(regB[23]), .QN(n463) );
  DFF_X1 regB_reg_22_ ( .D(n322), .CK(clk), .Q(MB[22]), .QN(n464) );
  DFF_X1 regB_reg_21_ ( .D(n321), .CK(clk), .Q(MB[21]), .QN(n465) );
  DFF_X1 regB_reg_20_ ( .D(n320), .CK(clk), .Q(MB[20]), .QN(n466) );
  DFF_X1 regB_reg_19_ ( .D(n319), .CK(clk), .Q(MB[19]), .QN(n467) );
  DFF_X1 regB_reg_18_ ( .D(n318), .CK(clk), .Q(MB[18]), .QN(n468) );
  DFF_X1 regB_reg_17_ ( .D(n317), .CK(clk), .Q(MB[17]), .QN(n469) );
  DFF_X1 regB_reg_16_ ( .D(n316), .CK(clk), .Q(MB[16]), .QN(n470) );
  DFF_X1 regB_reg_15_ ( .D(n315), .CK(clk), .Q(MB[15]), .QN(n471) );
  DFF_X1 regB_reg_14_ ( .D(n314), .CK(clk), .Q(MB[14]), .QN(n472) );
  DFF_X1 regB_reg_13_ ( .D(n313), .CK(clk), .Q(MB[13]), .QN(n473) );
  DFF_X1 regB_reg_12_ ( .D(n312), .CK(clk), .Q(MB[12]), .QN(n474) );
  DFF_X1 regB_reg_11_ ( .D(n311), .CK(clk), .Q(MB[11]), .QN(n475) );
  DFF_X1 regB_reg_10_ ( .D(n310), .CK(clk), .Q(MB[10]), .QN(n476) );
  DFF_X1 regB_reg_9_ ( .D(n309), .CK(clk), .Q(MB[9]), .QN(n477) );
  DFF_X1 regB_reg_8_ ( .D(n308), .CK(clk), .Q(MB[8]), .QN(n478) );
  DFF_X1 regB_reg_7_ ( .D(n307), .CK(clk), .Q(MB[7]), .QN(n479) );
  DFF_X1 regB_reg_6_ ( .D(n306), .CK(clk), .Q(MB[6]), .QN(n480) );
  DFF_X1 regB_reg_5_ ( .D(n305), .CK(clk), .Q(MB[5]), .QN(n481) );
  DFF_X1 regB_reg_4_ ( .D(n304), .CK(clk), .Q(MB[4]), .QN(n482) );
  DFF_X1 regB_reg_3_ ( .D(n303), .CK(clk), .Q(MB[3]), .QN(n483) );
  DFF_X1 regB_reg_2_ ( .D(n302), .CK(clk), .Q(MB[2]), .QN(n484) );
  DFF_X1 regB_reg_1_ ( .D(n301), .CK(clk), .Q(MB[1]), .QN(n485) );
  DFF_X1 regB_reg_0_ ( .D(n300), .CK(clk), .Q(MB[0]), .QN(n486) );
  DFF_X1 regA_reg_31_ ( .D(n299), .CK(clk), .Q(n200), .QN(n487) );
  DFF_X1 regA_reg_30_ ( .D(n298), .CK(clk), .Q(regA[30]), .QN(n488) );
  DFF_X1 regA_reg_29_ ( .D(n297), .CK(clk), .Q(regA[29]), .QN(n489) );
  DFF_X1 regA_reg_28_ ( .D(n296), .CK(clk), .Q(regA[28]), .QN(n490) );
  DFF_X1 regA_reg_27_ ( .D(n295), .CK(clk), .Q(regA[27]), .QN(n491) );
  DFF_X1 regA_reg_26_ ( .D(n294), .CK(clk), .Q(regA[26]), .QN(n492) );
  DFF_X1 regA_reg_25_ ( .D(n293), .CK(clk), .Q(regA[25]), .QN(n493) );
  DFF_X1 regA_reg_24_ ( .D(n292), .CK(clk), .Q(regA[24]), .QN(n494) );
  DFF_X1 regA_reg_23_ ( .D(n291), .CK(clk), .Q(regA[23]), .QN(n495) );
  DFF_X1 regA_reg_22_ ( .D(n290), .CK(clk), .Q(MA[22]), .QN(n496) );
  DFF_X1 regA_reg_21_ ( .D(n289), .CK(clk), .Q(MA[21]), .QN(n497) );
  DFF_X1 regA_reg_20_ ( .D(n288), .CK(clk), .Q(MA[20]), .QN(n498) );
  DFF_X1 regA_reg_19_ ( .D(n287), .CK(clk), .Q(MA[19]), .QN(n499) );
  DFF_X1 regA_reg_18_ ( .D(n286), .CK(clk), .Q(MA[18]), .QN(n500) );
  DFF_X1 regA_reg_17_ ( .D(n285), .CK(clk), .Q(MA[17]), .QN(n501) );
  DFF_X1 regA_reg_16_ ( .D(n284), .CK(clk), .Q(MA[16]), .QN(n502) );
  DFF_X1 regA_reg_15_ ( .D(n283), .CK(clk), .Q(MA[15]), .QN(n503) );
  DFF_X1 regA_reg_14_ ( .D(n282), .CK(clk), .Q(MA[14]), .QN(n504) );
  DFF_X1 regA_reg_13_ ( .D(n281), .CK(clk), .Q(MA[13]), .QN(n505) );
  DFF_X1 regA_reg_12_ ( .D(n280), .CK(clk), .Q(MA[12]), .QN(n506) );
  DFF_X1 regA_reg_11_ ( .D(n279), .CK(clk), .Q(MA[11]), .QN(n507) );
  DFF_X1 regA_reg_10_ ( .D(n278), .CK(clk), .Q(MA[10]), .QN(n508) );
  DFF_X1 regA_reg_9_ ( .D(n277), .CK(clk), .Q(MA[9]), .QN(n509) );
  DFF_X1 regA_reg_8_ ( .D(n276), .CK(clk), .Q(MA[8]), .QN(n510) );
  DFF_X1 regA_reg_7_ ( .D(n275), .CK(clk), .Q(MA[7]), .QN(n511) );
  DFF_X1 regA_reg_6_ ( .D(n274), .CK(clk), .Q(MA[6]), .QN(n512) );
  DFF_X1 regA_reg_5_ ( .D(n273), .CK(clk), .Q(MA[5]), .QN(n513) );
  DFF_X1 regA_reg_4_ ( .D(n272), .CK(clk), .Q(MA[4]), .QN(n514) );
  DFF_X1 regA_reg_3_ ( .D(n271), .CK(clk), .Q(MA[3]), .QN(n515) );
  DFF_X1 regA_reg_2_ ( .D(n270), .CK(clk), .Q(MA[2]), .QN(n516) );
  DFF_X1 regA_reg_1_ ( .D(n269), .CK(clk), .Q(MA[1]), .QN(n517) );
  DFF_X1 regA_reg_0_ ( .D(n268), .CK(clk), .Q(MA[0]), .QN(n518) );
  XNOR2_X1 U294 ( .A(add_0_root_sub_1_root_add_24_2_A_6_), .B(n344), .ZN(n332)
         );
  XNOR2_X1 U295 ( .A(add_0_root_sub_1_root_add_24_2_A_2_), .B(
        add_0_root_sub_1_root_add_24_2_carry_2_), .ZN(n333) );
  XNOR2_X1 U296 ( .A(add_0_root_sub_1_root_add_24_2_A_3_), .B(n341), .ZN(n334)
         );
  XNOR2_X1 U297 ( .A(add_0_root_sub_1_root_add_24_2_A_4_), .B(n342), .ZN(n335)
         );
  XNOR2_X1 U298 ( .A(add_0_root_sub_1_root_add_24_2_A_5_), .B(n343), .ZN(n336)
         );
  XNOR2_X1 U299 ( .A(N80), .B(add_0_root_sub_1_root_add_24_2_A_0_), .ZN(n337)
         );
  XOR2_X1 U300 ( .A(add_0_root_sub_1_root_add_24_2_A_8_), .B(n338), .Z(n346)
         );
  NAND2_X1 U301 ( .A1(n347), .A2(n348), .ZN(n338) );
  XOR2_X1 U302 ( .A(add_0_root_sub_1_root_add_24_2_A_7_), .B(n345), .Z(n339)
         );
  INV_X1 U303 ( .A(mantissasProduct[44]), .ZN(n369) );
  INV_X1 U304 ( .A(mantissasProduct[43]), .ZN(n370) );
  INV_X1 U305 ( .A(mantissasProduct[30]), .ZN(n383) );
  INV_X1 U306 ( .A(mantissasProduct[32]), .ZN(n381) );
  INV_X1 U307 ( .A(mantissasProduct[34]), .ZN(n379) );
  INV_X1 U308 ( .A(mantissasProduct[36]), .ZN(n377) );
  INV_X1 U309 ( .A(mantissasProduct[38]), .ZN(n375) );
  INV_X1 U310 ( .A(mantissasProduct[40]), .ZN(n373) );
  INV_X1 U311 ( .A(mantissasProduct[42]), .ZN(n371) );
  INV_X1 U312 ( .A(mantissasProduct[28]), .ZN(n385) );
  INV_X1 U313 ( .A(mantissasProduct[27]), .ZN(n386) );
  INV_X1 U314 ( .A(mantissasProduct[29]), .ZN(n384) );
  INV_X1 U315 ( .A(mantissasProduct[31]), .ZN(n382) );
  INV_X1 U316 ( .A(mantissasProduct[33]), .ZN(n380) );
  INV_X1 U317 ( .A(mantissasProduct[35]), .ZN(n378) );
  INV_X1 U318 ( .A(mantissasProduct[39]), .ZN(n374) );
  INV_X1 U319 ( .A(mantissasProduct[41]), .ZN(n372) );
  INV_X1 U320 ( .A(mantissasProduct[37]), .ZN(n376) );
  INV_X1 U321 ( .A(mantissasProduct[25]), .ZN(n388) );
  INV_X1 U322 ( .A(mantissasProduct[26]), .ZN(n387) );
  BUF_X1 U323 ( .A(n349), .Z(n351) );
  BUF_X1 U324 ( .A(n349), .Z(n352) );
  BUF_X1 U325 ( .A(n349), .Z(n353) );
  BUF_X1 U326 ( .A(n350), .Z(n354) );
  BUF_X1 U327 ( .A(n350), .Z(n355) );
  INV_X1 U328 ( .A(n142), .ZN(n367) );
  INV_X1 U329 ( .A(n143), .ZN(n366) );
  INV_X1 U330 ( .A(n345), .ZN(n348) );
  NOR2_X1 U331 ( .A1(N80), .A2(n9), .ZN(n143) );
  AND2_X1 U332 ( .A1(N80), .A2(add_0_root_sub_1_root_add_24_2_A_0_), .ZN(n340)
         );
  AND2_X1 U333 ( .A1(add_0_root_sub_1_root_add_24_2_A_2_), .A2(
        add_0_root_sub_1_root_add_24_2_carry_2_), .ZN(n341) );
  AND2_X1 U334 ( .A1(add_0_root_sub_1_root_add_24_2_A_3_), .A2(n341), .ZN(n342) );
  AND2_X1 U335 ( .A1(add_0_root_sub_1_root_add_24_2_A_4_), .A2(n342), .ZN(n343) );
  AND2_X1 U336 ( .A1(add_0_root_sub_1_root_add_24_2_A_5_), .A2(n343), .ZN(n344) );
  AND2_X1 U337 ( .A1(add_0_root_sub_1_root_add_24_2_A_6_), .A2(n344), .ZN(n345) );
  INV_X1 U338 ( .A(add_0_root_sub_1_root_add_24_2_A_7_), .ZN(n347) );
  NAND3_X1 U339 ( .A1(n468), .A2(n467), .A3(n469), .ZN(n194) );
  NAND2_X1 U340 ( .A1(n364), .A2(n390), .ZN(n11) );
  OAI22_X1 U341 ( .A1(n364), .A2(n204), .B1(n9), .B2(n332), .ZN(n265) );
  OAI22_X1 U342 ( .A1(n364), .A2(n203), .B1(n9), .B2(n339), .ZN(n266) );
  OAI22_X1 U343 ( .A1(n364), .A2(n210), .B1(n9), .B2(n337), .ZN(n259) );
  OAI22_X1 U344 ( .A1(n364), .A2(n209), .B1(n9), .B2(n365), .ZN(n260) );
  INV_X1 U345 ( .A(N27), .ZN(n365) );
  OAI22_X1 U346 ( .A1(n363), .A2(n208), .B1(n9), .B2(n333), .ZN(n261) );
  OAI22_X1 U347 ( .A1(n364), .A2(n207), .B1(n9), .B2(n334), .ZN(n262) );
  OAI22_X1 U348 ( .A1(n364), .A2(n206), .B1(n9), .B2(n335), .ZN(n263) );
  OAI22_X1 U349 ( .A1(n363), .A2(n205), .B1(n9), .B2(n336), .ZN(n264) );
  OAI222_X1 U350 ( .A1(n366), .A2(n388), .B1(n367), .B2(n389), .C1(n358), .C2(
        n232), .ZN(n237) );
  INV_X1 U351 ( .A(mantissasProduct[24]), .ZN(n389) );
  OAI222_X1 U352 ( .A1(n366), .A2(n387), .B1(n367), .B2(n388), .C1(n358), .C2(
        n231), .ZN(n238) );
  OAI222_X1 U353 ( .A1(n366), .A2(n386), .B1(n367), .B2(n387), .C1(n358), .C2(
        n230), .ZN(n239) );
  OAI222_X1 U354 ( .A1(n366), .A2(n385), .B1(n367), .B2(n386), .C1(n358), .C2(
        n229), .ZN(n240) );
  OAI222_X1 U355 ( .A1(n366), .A2(n384), .B1(n367), .B2(n385), .C1(n358), .C2(
        n228), .ZN(n241) );
  OAI222_X1 U356 ( .A1(n366), .A2(n383), .B1(n367), .B2(n384), .C1(n357), .C2(
        n227), .ZN(n242) );
  OAI222_X1 U357 ( .A1(n366), .A2(n382), .B1(n367), .B2(n383), .C1(n358), .C2(
        n226), .ZN(n243) );
  OAI222_X1 U358 ( .A1(n366), .A2(n381), .B1(n367), .B2(n382), .C1(n357), .C2(
        n225), .ZN(n244) );
  OAI222_X1 U359 ( .A1(n366), .A2(n380), .B1(n367), .B2(n381), .C1(n357), .C2(
        n224), .ZN(n245) );
  OAI222_X1 U360 ( .A1(n366), .A2(n379), .B1(n367), .B2(n380), .C1(n358), .C2(
        n223), .ZN(n246) );
  OAI222_X1 U361 ( .A1(n366), .A2(n378), .B1(n367), .B2(n379), .C1(n357), .C2(
        n222), .ZN(n247) );
  OAI222_X1 U362 ( .A1(n366), .A2(n377), .B1(n367), .B2(n378), .C1(n358), .C2(
        n221), .ZN(n248) );
  OAI222_X1 U363 ( .A1(n366), .A2(n376), .B1(n367), .B2(n377), .C1(n357), .C2(
        n220), .ZN(n249) );
  OAI222_X1 U364 ( .A1(n366), .A2(n375), .B1(n367), .B2(n376), .C1(n358), .C2(
        n219), .ZN(n250) );
  OAI222_X1 U365 ( .A1(n366), .A2(n374), .B1(n367), .B2(n375), .C1(n357), .C2(
        n218), .ZN(n251) );
  OAI222_X1 U366 ( .A1(n366), .A2(n373), .B1(n367), .B2(n374), .C1(n357), .C2(
        n217), .ZN(n252) );
  OAI222_X1 U367 ( .A1(n366), .A2(n372), .B1(n367), .B2(n373), .C1(n357), .C2(
        n216), .ZN(n253) );
  OAI222_X1 U368 ( .A1(n366), .A2(n371), .B1(n367), .B2(n372), .C1(n357), .C2(
        n215), .ZN(n254) );
  OAI222_X1 U369 ( .A1(n366), .A2(n370), .B1(n367), .B2(n371), .C1(n357), .C2(
        n214), .ZN(n255) );
  OAI222_X1 U370 ( .A1(n366), .A2(n369), .B1(n367), .B2(n370), .C1(n357), .C2(
        n213), .ZN(n256) );
  OAI222_X1 U371 ( .A1(n366), .A2(n368), .B1(n367), .B2(n369), .C1(n357), .C2(
        n212), .ZN(n257) );
  INV_X1 U372 ( .A(mantissasProduct[45]), .ZN(n368) );
  OAI21_X1 U373 ( .B1(n364), .B2(n233), .A(n141), .ZN(n236) );
  AOI22_X1 U374 ( .A1(mantissasProduct[23]), .A2(n142), .B1(
        mantissasProduct[24]), .B2(n143), .ZN(n141) );
  NOR4_X1 U375 ( .A1(regB[30]), .A2(regB[29]), .A3(regB[28]), .A4(regB[27]), 
        .ZN(n197) );
  OAI21_X1 U376 ( .B1(n364), .B2(n211), .A(n168), .ZN(n258) );
  AOI22_X1 U377 ( .A1(mantissasProduct[45]), .A2(n142), .B1(
        mantissasProduct[46]), .B2(n143), .ZN(n168) );
  NAND2_X1 U378 ( .A1(n198), .A2(n199), .ZN(MA[23]) );
  NOR4_X1 U379 ( .A1(regA[30]), .A2(regA[29]), .A3(regA[28]), .A4(regA[27]), 
        .ZN(n199) );
  NOR4_X1 U380 ( .A1(regA[26]), .A2(regA[25]), .A3(regA[24]), .A4(regA[23]), 
        .ZN(n198) );
  NAND4_X1 U381 ( .A1(n364), .A2(n178), .A3(n179), .A4(n390), .ZN(n9) );
  NAND4_X1 U382 ( .A1(n188), .A2(n189), .A3(n190), .A4(n191), .ZN(n178) );
  NAND4_X1 U383 ( .A1(n180), .A2(n181), .A3(n182), .A4(n183), .ZN(n179) );
  NOR4_X1 U384 ( .A1(n194), .A2(MB[14]), .A3(MB[16]), .A4(MB[15]), .ZN(n189)
         );
  NOR4_X1 U385 ( .A1(n184), .A2(MA[4]), .A3(MA[6]), .A4(MA[5]), .ZN(n183) );
  NAND4_X1 U386 ( .A1(n511), .A2(n510), .A3(n509), .A4(n487), .ZN(n184) );
  NOR4_X1 U387 ( .A1(n185), .A2(MA[1]), .A3(MA[21]), .A4(MA[20]), .ZN(n182) );
  NAND3_X1 U388 ( .A1(n516), .A2(n515), .A3(n496), .ZN(n185) );
  NOR4_X1 U389 ( .A1(n193), .A2(MB[1]), .A3(MB[21]), .A4(MB[20]), .ZN(n190) );
  NAND3_X1 U390 ( .A1(n484), .A2(n483), .A3(n464), .ZN(n193) );
  NOR4_X1 U391 ( .A1(n187), .A2(MA[23]), .A3(MA[10]), .A4(MA[0]), .ZN(n180) );
  NAND3_X1 U392 ( .A1(n506), .A2(n505), .A3(n507), .ZN(n187) );
  NOR4_X1 U393 ( .A1(n195), .A2(MB[23]), .A3(MB[10]), .A4(MB[0]), .ZN(n188) );
  NAND3_X1 U394 ( .A1(n474), .A2(n473), .A3(n475), .ZN(n195) );
  BUF_X1 U395 ( .A(enable), .Z(n359) );
  BUF_X1 U396 ( .A(enable), .Z(n360) );
  BUF_X1 U397 ( .A(enable), .Z(n361) );
  BUF_X1 U398 ( .A(enable), .Z(n362) );
  BUF_X1 U399 ( .A(enable), .Z(n357) );
  BUF_X1 U400 ( .A(enable), .Z(n358) );
  BUF_X1 U401 ( .A(enable), .Z(n363) );
  OAI22_X1 U402 ( .A1(n361), .A2(n202), .B1(n8), .B2(n9), .ZN(n267) );
  XNOR2_X1 U403 ( .A(n201), .B(n200), .ZN(n8) );
  BUF_X1 U404 ( .A(enable), .Z(n364) );
  INV_X1 U405 ( .A(B[23]), .ZN(n431) );
  INV_X1 U406 ( .A(B[27]), .ZN(n427) );
  NOR4_X1 U407 ( .A1(n192), .A2(MB[4]), .A3(MB[6]), .A4(MB[5]), .ZN(n191) );
  NAND4_X1 U408 ( .A1(n479), .A2(n478), .A3(n477), .A4(n455), .ZN(n192) );
  OAI22_X1 U409 ( .A1(n363), .A2(n458), .B1(n356), .B2(n426), .ZN(n328) );
  INV_X1 U410 ( .A(B[28]), .ZN(n426) );
  OAI22_X1 U411 ( .A1(n363), .A2(n457), .B1(n356), .B2(n425), .ZN(n329) );
  INV_X1 U412 ( .A(B[29]), .ZN(n425) );
  OAI22_X1 U413 ( .A1(n363), .A2(n456), .B1(n356), .B2(n424), .ZN(n330) );
  INV_X1 U414 ( .A(B[30]), .ZN(n424) );
  OAI22_X1 U415 ( .A1(n363), .A2(n455), .B1(n356), .B2(n423), .ZN(n331) );
  INV_X1 U416 ( .A(B[31]), .ZN(n423) );
  OAI22_X1 U417 ( .A1(n359), .A2(n518), .B1(n351), .B2(n422), .ZN(n268) );
  INV_X1 U418 ( .A(A[0]), .ZN(n422) );
  OAI22_X1 U419 ( .A1(n358), .A2(n517), .B1(n351), .B2(n421), .ZN(n269) );
  INV_X1 U420 ( .A(A[1]), .ZN(n421) );
  OAI22_X1 U421 ( .A1(n359), .A2(n516), .B1(n351), .B2(n420), .ZN(n270) );
  INV_X1 U422 ( .A(A[2]), .ZN(n420) );
  OAI22_X1 U423 ( .A1(n359), .A2(n515), .B1(n351), .B2(n419), .ZN(n271) );
  INV_X1 U424 ( .A(A[3]), .ZN(n419) );
  OAI22_X1 U425 ( .A1(n359), .A2(n514), .B1(n351), .B2(n418), .ZN(n272) );
  INV_X1 U426 ( .A(A[4]), .ZN(n418) );
  OAI22_X1 U427 ( .A1(n358), .A2(n513), .B1(n351), .B2(n417), .ZN(n273) );
  INV_X1 U428 ( .A(A[5]), .ZN(n417) );
  OAI22_X1 U429 ( .A1(n359), .A2(n512), .B1(n351), .B2(n416), .ZN(n274) );
  INV_X1 U430 ( .A(A[6]), .ZN(n416) );
  OAI22_X1 U431 ( .A1(n358), .A2(n511), .B1(n351), .B2(n415), .ZN(n275) );
  INV_X1 U432 ( .A(A[7]), .ZN(n415) );
  OAI22_X1 U433 ( .A1(n359), .A2(n510), .B1(n351), .B2(n414), .ZN(n276) );
  INV_X1 U434 ( .A(A[8]), .ZN(n414) );
  OAI22_X1 U435 ( .A1(n359), .A2(n509), .B1(n351), .B2(n413), .ZN(n277) );
  INV_X1 U436 ( .A(A[9]), .ZN(n413) );
  OAI22_X1 U437 ( .A1(n359), .A2(n508), .B1(n351), .B2(n412), .ZN(n278) );
  INV_X1 U438 ( .A(A[10]), .ZN(n412) );
  OAI22_X1 U439 ( .A1(n359), .A2(n507), .B1(n351), .B2(n411), .ZN(n279) );
  INV_X1 U440 ( .A(A[11]), .ZN(n411) );
  OAI22_X1 U441 ( .A1(n359), .A2(n506), .B1(n352), .B2(n410), .ZN(n280) );
  INV_X1 U442 ( .A(A[12]), .ZN(n410) );
  OAI22_X1 U443 ( .A1(n359), .A2(n505), .B1(n352), .B2(n409), .ZN(n281) );
  INV_X1 U444 ( .A(A[13]), .ZN(n409) );
  OAI22_X1 U445 ( .A1(n359), .A2(n504), .B1(n352), .B2(n408), .ZN(n282) );
  INV_X1 U446 ( .A(A[14]), .ZN(n408) );
  OAI22_X1 U447 ( .A1(n359), .A2(n503), .B1(n352), .B2(n407), .ZN(n283) );
  INV_X1 U448 ( .A(A[15]), .ZN(n407) );
  OAI22_X1 U449 ( .A1(n360), .A2(n502), .B1(n352), .B2(n406), .ZN(n284) );
  INV_X1 U450 ( .A(A[16]), .ZN(n406) );
  OAI22_X1 U451 ( .A1(n360), .A2(n501), .B1(n352), .B2(n405), .ZN(n285) );
  INV_X1 U452 ( .A(A[17]), .ZN(n405) );
  OAI22_X1 U453 ( .A1(n360), .A2(n500), .B1(n352), .B2(n404), .ZN(n286) );
  INV_X1 U454 ( .A(A[18]), .ZN(n404) );
  OAI22_X1 U455 ( .A1(n360), .A2(n499), .B1(n352), .B2(n403), .ZN(n287) );
  INV_X1 U456 ( .A(A[19]), .ZN(n403) );
  OAI22_X1 U457 ( .A1(n360), .A2(n498), .B1(n352), .B2(n402), .ZN(n288) );
  INV_X1 U458 ( .A(A[20]), .ZN(n402) );
  OAI22_X1 U459 ( .A1(n360), .A2(n497), .B1(n352), .B2(n401), .ZN(n289) );
  INV_X1 U460 ( .A(A[21]), .ZN(n401) );
  OAI22_X1 U461 ( .A1(n360), .A2(n496), .B1(n352), .B2(n400), .ZN(n290) );
  INV_X1 U462 ( .A(A[22]), .ZN(n400) );
  OAI22_X1 U463 ( .A1(n360), .A2(n495), .B1(n352), .B2(n399), .ZN(n291) );
  INV_X1 U464 ( .A(A[23]), .ZN(n399) );
  OAI22_X1 U465 ( .A1(n360), .A2(n494), .B1(n353), .B2(n398), .ZN(n292) );
  INV_X1 U466 ( .A(A[24]), .ZN(n398) );
  OAI22_X1 U467 ( .A1(n360), .A2(n493), .B1(n353), .B2(n397), .ZN(n293) );
  INV_X1 U468 ( .A(A[25]), .ZN(n397) );
  OAI22_X1 U469 ( .A1(n360), .A2(n492), .B1(n353), .B2(n396), .ZN(n294) );
  INV_X1 U470 ( .A(A[26]), .ZN(n396) );
  OAI22_X1 U471 ( .A1(n360), .A2(n491), .B1(n353), .B2(n395), .ZN(n295) );
  INV_X1 U472 ( .A(A[27]), .ZN(n395) );
  OAI22_X1 U473 ( .A1(n360), .A2(n490), .B1(n353), .B2(n394), .ZN(n296) );
  INV_X1 U474 ( .A(A[28]), .ZN(n394) );
  OAI22_X1 U475 ( .A1(n361), .A2(n489), .B1(n353), .B2(n393), .ZN(n297) );
  INV_X1 U476 ( .A(A[29]), .ZN(n393) );
  OAI22_X1 U477 ( .A1(n361), .A2(n488), .B1(n353), .B2(n392), .ZN(n298) );
  INV_X1 U478 ( .A(A[30]), .ZN(n392) );
  OAI22_X1 U479 ( .A1(n361), .A2(n487), .B1(n353), .B2(n391), .ZN(n299) );
  INV_X1 U480 ( .A(A[31]), .ZN(n391) );
  OAI22_X1 U481 ( .A1(n361), .A2(n486), .B1(n353), .B2(n454), .ZN(n300) );
  INV_X1 U482 ( .A(B[0]), .ZN(n454) );
  OAI22_X1 U483 ( .A1(n361), .A2(n485), .B1(n353), .B2(n453), .ZN(n301) );
  INV_X1 U484 ( .A(B[1]), .ZN(n453) );
  OAI22_X1 U485 ( .A1(n361), .A2(n484), .B1(n353), .B2(n452), .ZN(n302) );
  INV_X1 U486 ( .A(B[2]), .ZN(n452) );
  OAI22_X1 U487 ( .A1(n361), .A2(n483), .B1(n353), .B2(n451), .ZN(n303) );
  INV_X1 U488 ( .A(B[3]), .ZN(n451) );
  OAI22_X1 U489 ( .A1(n361), .A2(n482), .B1(n354), .B2(n450), .ZN(n304) );
  INV_X1 U490 ( .A(B[4]), .ZN(n450) );
  OAI22_X1 U491 ( .A1(n361), .A2(n481), .B1(n354), .B2(n449), .ZN(n305) );
  INV_X1 U492 ( .A(B[5]), .ZN(n449) );
  OAI22_X1 U493 ( .A1(n361), .A2(n480), .B1(n354), .B2(n448), .ZN(n306) );
  INV_X1 U494 ( .A(B[6]), .ZN(n448) );
  OAI22_X1 U495 ( .A1(n361), .A2(n479), .B1(n354), .B2(n447), .ZN(n307) );
  INV_X1 U496 ( .A(B[7]), .ZN(n447) );
  OAI22_X1 U497 ( .A1(n361), .A2(n478), .B1(n354), .B2(n446), .ZN(n308) );
  INV_X1 U498 ( .A(B[8]), .ZN(n446) );
  OAI22_X1 U499 ( .A1(n362), .A2(n477), .B1(n354), .B2(n445), .ZN(n309) );
  INV_X1 U500 ( .A(B[9]), .ZN(n445) );
  OAI22_X1 U501 ( .A1(n362), .A2(n476), .B1(n354), .B2(n444), .ZN(n310) );
  INV_X1 U502 ( .A(B[10]), .ZN(n444) );
  OAI22_X1 U503 ( .A1(n362), .A2(n475), .B1(n354), .B2(n443), .ZN(n311) );
  INV_X1 U504 ( .A(B[11]), .ZN(n443) );
  OAI22_X1 U505 ( .A1(n362), .A2(n474), .B1(n354), .B2(n442), .ZN(n312) );
  INV_X1 U506 ( .A(B[12]), .ZN(n442) );
  OAI22_X1 U507 ( .A1(n362), .A2(n473), .B1(n354), .B2(n441), .ZN(n313) );
  INV_X1 U508 ( .A(B[13]), .ZN(n441) );
  OAI22_X1 U509 ( .A1(n362), .A2(n472), .B1(n354), .B2(n440), .ZN(n314) );
  INV_X1 U510 ( .A(B[14]), .ZN(n440) );
  OAI22_X1 U511 ( .A1(n362), .A2(n471), .B1(n354), .B2(n439), .ZN(n315) );
  INV_X1 U512 ( .A(B[15]), .ZN(n439) );
  OAI22_X1 U513 ( .A1(n362), .A2(n470), .B1(n355), .B2(n438), .ZN(n316) );
  INV_X1 U514 ( .A(B[16]), .ZN(n438) );
  OAI22_X1 U515 ( .A1(n362), .A2(n469), .B1(n355), .B2(n437), .ZN(n317) );
  INV_X1 U516 ( .A(B[17]), .ZN(n437) );
  OAI22_X1 U517 ( .A1(n362), .A2(n468), .B1(n355), .B2(n436), .ZN(n318) );
  INV_X1 U518 ( .A(B[18]), .ZN(n436) );
  OAI22_X1 U519 ( .A1(n362), .A2(n467), .B1(n355), .B2(n435), .ZN(n319) );
  INV_X1 U520 ( .A(B[19]), .ZN(n435) );
  OAI22_X1 U521 ( .A1(n362), .A2(n466), .B1(n355), .B2(n434), .ZN(n320) );
  INV_X1 U522 ( .A(B[20]), .ZN(n434) );
  OAI22_X1 U523 ( .A1(n362), .A2(n465), .B1(n355), .B2(n433), .ZN(n321) );
  INV_X1 U524 ( .A(B[21]), .ZN(n433) );
  OAI22_X1 U525 ( .A1(n363), .A2(n464), .B1(n355), .B2(n432), .ZN(n322) );
  INV_X1 U526 ( .A(B[22]), .ZN(n432) );
  OAI22_X1 U527 ( .A1(n363), .A2(n462), .B1(n355), .B2(n430), .ZN(n324) );
  INV_X1 U528 ( .A(B[24]), .ZN(n430) );
  OAI22_X1 U529 ( .A1(n363), .A2(n461), .B1(n355), .B2(n429), .ZN(n325) );
  INV_X1 U530 ( .A(B[25]), .ZN(n429) );
  OAI22_X1 U531 ( .A1(n363), .A2(n460), .B1(n355), .B2(n428), .ZN(n326) );
  INV_X1 U532 ( .A(B[26]), .ZN(n428) );
  NOR4_X1 U533 ( .A1(n186), .A2(MA[14]), .A3(MA[16]), .A4(MA[15]), .ZN(n181)
         );
  NAND3_X1 U534 ( .A1(n500), .A2(n499), .A3(n501), .ZN(n186) );
  INV_X1 U535 ( .A(reset), .ZN(n390) );
  OAI22_X1 U536 ( .A1(n363), .A2(n463), .B1(n355), .B2(n431), .ZN(n323) );
  OAI22_X1 U537 ( .A1(n363), .A2(n459), .B1(n355), .B2(n427), .ZN(n327) );
  NOR4_X1 U538 ( .A1(regB[26]), .A2(regB[25]), .A3(regB[24]), .A4(regB[23]), 
        .ZN(n196) );
  NOR2_X1 U539 ( .A1(n9), .A2(N90), .ZN(n142) );
  NAND2_X1 U540 ( .A1(n196), .A2(n197), .ZN(MB[23]) );
  INV_X1 U541 ( .A(N90), .ZN(N80) );
  OAI22_X1 U542 ( .A1(n363), .A2(n234), .B1(n9), .B2(n346), .ZN(n235) );
  BUF_X1 U543 ( .A(n11), .Z(n349) );
  BUF_X1 U544 ( .A(n11), .Z(n350) );
  BUF_X1 U545 ( .A(n350), .Z(n356) );
endmodule

