
module fpAdder_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25;
  wire   [23:1] carry;

  FA_X1 U2_23 ( .A(A[23]), .B(n18), .CI(carry[23]), .S(DIFF[23]) );
  FA_X1 U2_22 ( .A(A[22]), .B(n17), .CI(carry[22]), .CO(carry[23]), .S(
        DIFF[22]) );
  FA_X1 U2_21 ( .A(A[21]), .B(n16), .CI(carry[21]), .CO(carry[22]), .S(
        DIFF[21]) );
  FA_X1 U2_20 ( .A(A[20]), .B(n15), .CI(carry[20]), .CO(carry[21]), .S(
        DIFF[20]) );
  FA_X1 U2_19 ( .A(A[19]), .B(n24), .CI(carry[19]), .CO(carry[20]), .S(
        DIFF[19]) );
  FA_X1 U2_18 ( .A(A[18]), .B(n23), .CI(carry[18]), .CO(carry[19]), .S(
        DIFF[18]) );
  FA_X1 U2_17 ( .A(A[17]), .B(n22), .CI(carry[17]), .CO(carry[18]), .S(
        DIFF[17]) );
  FA_X1 U2_16 ( .A(A[16]), .B(n21), .CI(carry[16]), .CO(carry[17]), .S(
        DIFF[16]) );
  FA_X1 U2_15 ( .A(A[15]), .B(n14), .CI(carry[15]), .CO(carry[16]), .S(
        DIFF[15]) );
  FA_X1 U2_14 ( .A(A[14]), .B(n13), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  FA_X1 U2_13 ( .A(A[13]), .B(n12), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  FA_X1 U2_12 ( .A(A[12]), .B(n11), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  FA_X1 U2_11 ( .A(A[11]), .B(n10), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  FA_X1 U2_10 ( .A(A[10]), .B(n9), .CI(carry[10]), .CO(carry[11]), .S(DIFF[10]) );
  FA_X1 U2_9 ( .A(A[9]), .B(n20), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  FA_X1 U2_8 ( .A(A[8]), .B(n19), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8]) );
  FA_X1 U2_7 ( .A(A[7]), .B(n5), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7]) );
  FA_X1 U2_6 ( .A(A[6]), .B(n4), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  FA_X1 U2_5 ( .A(A[5]), .B(n3), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  FA_X1 U2_4 ( .A(A[4]), .B(n2), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  FA_X1 U2_3 ( .A(A[3]), .B(n6), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  FA_X1 U2_2 ( .A(A[2]), .B(n7), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  FA_X1 U2_1 ( .A(A[1]), .B(n8), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  INV_X1 U1 ( .A(B[23]), .ZN(n18) );
  XNOR2_X1 U2 ( .A(n25), .B(A[0]), .ZN(DIFF[0]) );
  INV_X1 U3 ( .A(B[0]), .ZN(n25) );
  INV_X1 U4 ( .A(B[1]), .ZN(n8) );
  NAND2_X1 U5 ( .A1(B[0]), .A2(n1), .ZN(carry[1]) );
  INV_X1 U6 ( .A(A[0]), .ZN(n1) );
  INV_X1 U7 ( .A(B[2]), .ZN(n7) );
  INV_X1 U8 ( .A(B[3]), .ZN(n6) );
  INV_X1 U9 ( .A(B[4]), .ZN(n2) );
  INV_X1 U10 ( .A(B[5]), .ZN(n3) );
  INV_X1 U11 ( .A(B[6]), .ZN(n4) );
  INV_X1 U12 ( .A(B[7]), .ZN(n5) );
  INV_X1 U13 ( .A(B[8]), .ZN(n19) );
  INV_X1 U14 ( .A(B[9]), .ZN(n20) );
  INV_X1 U15 ( .A(B[10]), .ZN(n9) );
  INV_X1 U16 ( .A(B[11]), .ZN(n10) );
  INV_X1 U17 ( .A(B[12]), .ZN(n11) );
  INV_X1 U18 ( .A(B[13]), .ZN(n12) );
  INV_X1 U19 ( .A(B[14]), .ZN(n13) );
  INV_X1 U20 ( .A(B[15]), .ZN(n14) );
  INV_X1 U21 ( .A(B[16]), .ZN(n21) );
  INV_X1 U22 ( .A(B[17]), .ZN(n22) );
  INV_X1 U23 ( .A(B[18]), .ZN(n23) );
  INV_X1 U24 ( .A(B[19]), .ZN(n24) );
  INV_X1 U25 ( .A(B[20]), .ZN(n15) );
  INV_X1 U26 ( .A(B[21]), .ZN(n16) );
  INV_X1 U27 ( .A(B[22]), .ZN(n17) );
endmodule


module fpAdder_DW01_sub_2 ( A, B, CI, DIFF, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25;
  wire   [23:1] carry;

  FA_X1 U2_23 ( .A(A[23]), .B(n18), .CI(carry[23]), .S(DIFF[23]) );
  FA_X1 U2_22 ( .A(A[22]), .B(n17), .CI(carry[22]), .CO(carry[23]), .S(
        DIFF[22]) );
  FA_X1 U2_21 ( .A(A[21]), .B(n16), .CI(carry[21]), .CO(carry[22]), .S(
        DIFF[21]) );
  FA_X1 U2_20 ( .A(A[20]), .B(n15), .CI(carry[20]), .CO(carry[21]), .S(
        DIFF[20]) );
  FA_X1 U2_19 ( .A(A[19]), .B(n24), .CI(carry[19]), .CO(carry[20]), .S(
        DIFF[19]) );
  FA_X1 U2_18 ( .A(A[18]), .B(n23), .CI(carry[18]), .CO(carry[19]), .S(
        DIFF[18]) );
  FA_X1 U2_17 ( .A(A[17]), .B(n22), .CI(carry[17]), .CO(carry[18]), .S(
        DIFF[17]) );
  FA_X1 U2_16 ( .A(A[16]), .B(n21), .CI(carry[16]), .CO(carry[17]), .S(
        DIFF[16]) );
  FA_X1 U2_15 ( .A(A[15]), .B(n14), .CI(carry[15]), .CO(carry[16]), .S(
        DIFF[15]) );
  FA_X1 U2_14 ( .A(A[14]), .B(n13), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  FA_X1 U2_13 ( .A(A[13]), .B(n12), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  FA_X1 U2_12 ( .A(A[12]), .B(n11), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  FA_X1 U2_11 ( .A(A[11]), .B(n10), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  FA_X1 U2_10 ( .A(A[10]), .B(n9), .CI(carry[10]), .CO(carry[11]), .S(DIFF[10]) );
  FA_X1 U2_9 ( .A(A[9]), .B(n20), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  FA_X1 U2_8 ( .A(A[8]), .B(n19), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8]) );
  FA_X1 U2_7 ( .A(A[7]), .B(n5), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7]) );
  FA_X1 U2_6 ( .A(A[6]), .B(n4), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  FA_X1 U2_5 ( .A(A[5]), .B(n3), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  FA_X1 U2_4 ( .A(A[4]), .B(n2), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  FA_X1 U2_3 ( .A(A[3]), .B(n6), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  FA_X1 U2_2 ( .A(A[2]), .B(n7), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  FA_X1 U2_1 ( .A(A[1]), .B(n8), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  INV_X1 U1 ( .A(B[23]), .ZN(n18) );
  XNOR2_X1 U2 ( .A(n25), .B(A[0]), .ZN(DIFF[0]) );
  INV_X1 U3 ( .A(B[0]), .ZN(n25) );
  INV_X1 U4 ( .A(B[1]), .ZN(n8) );
  NAND2_X1 U5 ( .A1(B[0]), .A2(n1), .ZN(carry[1]) );
  INV_X1 U6 ( .A(A[0]), .ZN(n1) );
  INV_X1 U7 ( .A(B[2]), .ZN(n7) );
  INV_X1 U8 ( .A(B[3]), .ZN(n6) );
  INV_X1 U9 ( .A(B[4]), .ZN(n2) );
  INV_X1 U10 ( .A(B[5]), .ZN(n3) );
  INV_X1 U11 ( .A(B[6]), .ZN(n4) );
  INV_X1 U12 ( .A(B[7]), .ZN(n5) );
  INV_X1 U13 ( .A(B[8]), .ZN(n19) );
  INV_X1 U14 ( .A(B[9]), .ZN(n20) );
  INV_X1 U15 ( .A(B[10]), .ZN(n9) );
  INV_X1 U16 ( .A(B[11]), .ZN(n10) );
  INV_X1 U17 ( .A(B[12]), .ZN(n11) );
  INV_X1 U18 ( .A(B[13]), .ZN(n12) );
  INV_X1 U19 ( .A(B[14]), .ZN(n13) );
  INV_X1 U20 ( .A(B[15]), .ZN(n14) );
  INV_X1 U21 ( .A(B[16]), .ZN(n21) );
  INV_X1 U22 ( .A(B[17]), .ZN(n22) );
  INV_X1 U23 ( .A(B[18]), .ZN(n23) );
  INV_X1 U24 ( .A(B[19]), .ZN(n24) );
  INV_X1 U25 ( .A(B[20]), .ZN(n15) );
  INV_X1 U26 ( .A(B[21]), .ZN(n16) );
  INV_X1 U27 ( .A(B[22]), .ZN(n17) );
endmodule


module fpAdder_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HA_X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  HA_X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  HA_X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  HA_X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  HA_X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  HA_X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  INV_X1 U1 ( .A(A[0]), .ZN(SUM[0]) );
  XOR2_X1 U2 ( .A(carry[7]), .B(A[7]), .Z(SUM[7]) );
endmodule


module fpAdder_DW01_add_0 ( A, B, CI, SUM, CO );
  input [24:0] A;
  input [24:0] B;
  output [24:0] SUM;
  input CI;
  output CO;
  wire   n2;
  wire   [23:2] carry;

  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(SUM[24]), .S(SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n2), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U2 ( .A1(B[0]), .A2(A[0]), .ZN(n2) );
endmodule


module fpAdder_DW_rash_0 ( A, DATA_TC, SH, SH_TC, B );
  input [23:0] A;
  input [7:0] SH;
  output [23:0] B;
  input DATA_TC, SH_TC;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144;

  NAND2_X1 U3 ( .A1(n100), .A2(n10), .ZN(n61) );
  INV_X1 U4 ( .A(n122), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n91), .A2(n11), .ZN(n58) );
  BUF_X1 U6 ( .A(n97), .Z(n7) );
  BUF_X1 U7 ( .A(n97), .Z(n8) );
  INV_X1 U8 ( .A(n137), .ZN(n12) );
  INV_X1 U9 ( .A(n64), .ZN(n9) );
  INV_X1 U10 ( .A(n69), .ZN(n25) );
  INV_X1 U11 ( .A(n79), .ZN(n28) );
  INV_X1 U12 ( .A(n74), .ZN(n20) );
  INV_X1 U13 ( .A(SH[2]), .ZN(n13) );
  INV_X1 U14 ( .A(SH[0]), .ZN(n35) );
  INV_X1 U15 ( .A(n83), .ZN(n14) );
  INV_X1 U16 ( .A(SH[7]), .ZN(n11) );
  INV_X1 U17 ( .A(n87), .ZN(n17) );
  INV_X1 U18 ( .A(n80), .ZN(n31) );
  INV_X1 U19 ( .A(n77), .ZN(n29) );
  INV_X1 U20 ( .A(n84), .ZN(n15) );
  INV_X1 U21 ( .A(n72), .ZN(n21) );
  INV_X1 U22 ( .A(n67), .ZN(n26) );
  INV_X1 U23 ( .A(n65), .ZN(n23) );
  INV_X1 U24 ( .A(n85), .ZN(n18) );
  INV_X1 U25 ( .A(n78), .ZN(n27) );
  INV_X1 U26 ( .A(n73), .ZN(n22) );
  INV_X1 U27 ( .A(n102), .ZN(n24) );
  INV_X1 U28 ( .A(n112), .ZN(n19) );
  INV_X1 U29 ( .A(n88), .ZN(n16) );
  INV_X1 U30 ( .A(n75), .ZN(n32) );
  INV_X1 U31 ( .A(n81), .ZN(n30) );
  INV_X1 U32 ( .A(n70), .ZN(n33) );
  INV_X1 U33 ( .A(A[23]), .ZN(n36) );
  INV_X1 U34 ( .A(A[2]), .ZN(n57) );
  INV_X1 U35 ( .A(n94), .ZN(n34) );
  INV_X1 U36 ( .A(A[22]), .ZN(n37) );
  INV_X1 U37 ( .A(A[21]), .ZN(n38) );
  INV_X1 U38 ( .A(A[19]), .ZN(n40) );
  INV_X1 U39 ( .A(A[20]), .ZN(n39) );
  INV_X1 U40 ( .A(A[11]), .ZN(n48) );
  INV_X1 U41 ( .A(A[12]), .ZN(n47) );
  INV_X1 U42 ( .A(A[18]), .ZN(n41) );
  INV_X1 U43 ( .A(A[3]), .ZN(n56) );
  INV_X1 U44 ( .A(A[14]), .ZN(n45) );
  INV_X1 U45 ( .A(A[10]), .ZN(n49) );
  INV_X1 U46 ( .A(A[6]), .ZN(n53) );
  INV_X1 U47 ( .A(A[15]), .ZN(n44) );
  INV_X1 U48 ( .A(A[7]), .ZN(n52) );
  INV_X1 U49 ( .A(A[16]), .ZN(n43) );
  INV_X1 U50 ( .A(A[8]), .ZN(n51) );
  INV_X1 U51 ( .A(A[4]), .ZN(n55) );
  INV_X1 U52 ( .A(A[13]), .ZN(n46) );
  INV_X1 U53 ( .A(A[5]), .ZN(n54) );
  INV_X1 U54 ( .A(A[17]), .ZN(n42) );
  INV_X1 U55 ( .A(A[9]), .ZN(n50) );
  NOR2_X1 U56 ( .A1(n35), .A2(SH[1]), .ZN(n1) );
  NOR2_X1 U57 ( .A1(n35), .A2(SH[1]), .ZN(n2) );
  NAND2_X1 U58 ( .A1(n35), .A2(SH[1]), .ZN(n3) );
  NAND2_X1 U59 ( .A1(n35), .A2(SH[1]), .ZN(n4) );
  NAND2_X1 U60 ( .A1(SH[0]), .A2(SH[1]), .ZN(n5) );
  NAND2_X1 U61 ( .A1(SH[0]), .A2(SH[1]), .ZN(n6) );
  OAI222_X1 U62 ( .A1(n31), .A2(n58), .B1(n59), .B2(n60), .C1(n27), .C2(n61), 
        .ZN(B[9]) );
  OAI222_X1 U63 ( .A1(n17), .A2(n58), .B1(n62), .B2(n60), .C1(n18), .C2(n61), 
        .ZN(B[8]) );
  OAI221_X1 U64 ( .B1(n33), .B2(n58), .C1(n24), .C2(n61), .A(n63), .ZN(B[7])
         );
  AOI222_X1 U65 ( .A1(n64), .A2(n65), .B1(n66), .B2(n67), .C1(n68), .C2(n25), 
        .ZN(n63) );
  OAI221_X1 U66 ( .B1(n32), .B2(n58), .C1(n19), .C2(n61), .A(n71), .ZN(B[6])
         );
  AOI222_X1 U67 ( .A1(n68), .A2(n20), .B1(n66), .B2(n72), .C1(n64), .C2(n73), 
        .ZN(n71) );
  OAI221_X1 U68 ( .B1(n30), .B2(n58), .C1(n31), .C2(n61), .A(n76), .ZN(B[5])
         );
  AOI222_X1 U69 ( .A1(n68), .A2(n28), .B1(n66), .B2(n77), .C1(n64), .C2(n78), 
        .ZN(n76) );
  OAI221_X1 U70 ( .B1(n16), .B2(n58), .C1(n17), .C2(n61), .A(n82), .ZN(B[4])
         );
  AOI222_X1 U71 ( .A1(n68), .A2(n83), .B1(n66), .B2(n84), .C1(n64), .C2(n85), 
        .ZN(n82) );
  NOR2_X1 U72 ( .A1(n60), .A2(n13), .ZN(n66) );
  NOR4_X1 U73 ( .A1(n12), .A2(SH[2]), .A3(n86), .A4(SH[7]), .ZN(n68) );
  AOI21_X1 U74 ( .B1(n89), .B2(n90), .A(SH[7]), .ZN(B[3]) );
  NAND2_X1 U75 ( .A1(n91), .A2(n92), .ZN(n90) );
  OAI221_X1 U76 ( .B1(n93), .B2(n53), .C1(n3), .C2(n54), .A(n95), .ZN(n92) );
  AOI22_X1 U77 ( .A1(A[4]), .A2(n2), .B1(A[3]), .B2(n7), .ZN(n95) );
  MUX2_X1 U78 ( .A(n98), .B(n99), .S(n86), .Z(n89) );
  AOI222_X1 U79 ( .A1(n100), .A2(n70), .B1(n101), .B2(n102), .C1(n103), .C2(
        n65), .ZN(n99) );
  OAI221_X1 U80 ( .B1(n6), .B2(n49), .C1(n94), .C2(n50), .A(n104), .ZN(n70) );
  AOI22_X1 U81 ( .A1(A[8]), .A2(n1), .B1(A[7]), .B2(n7), .ZN(n104) );
  OR2_X1 U82 ( .A1(n12), .A2(n105), .ZN(n98) );
  AOI21_X1 U83 ( .B1(n106), .B2(n107), .A(SH[7]), .ZN(B[2]) );
  NAND2_X1 U84 ( .A1(n91), .A2(n108), .ZN(n107) );
  OAI221_X1 U85 ( .B1(n5), .B2(n54), .C1(n4), .C2(n55), .A(n109), .ZN(n108) );
  AOI22_X1 U86 ( .A1(A[3]), .A2(n96), .B1(A[2]), .B2(n7), .ZN(n109) );
  MUX2_X1 U87 ( .A(n110), .B(n111), .S(n86), .Z(n106) );
  AOI222_X1 U88 ( .A1(n100), .A2(n75), .B1(n101), .B2(n112), .C1(n103), .C2(
        n73), .ZN(n111) );
  OAI221_X1 U89 ( .B1(n93), .B2(n50), .C1(n3), .C2(n51), .A(n113), .ZN(n75) );
  AOI22_X1 U90 ( .A1(A[7]), .A2(n2), .B1(A[6]), .B2(n7), .ZN(n113) );
  NOR2_X1 U91 ( .A1(n58), .A2(n69), .ZN(B[23]) );
  NOR2_X1 U92 ( .A1(n74), .A2(n58), .ZN(B[22]) );
  NOR2_X1 U93 ( .A1(n79), .A2(n58), .ZN(B[21]) );
  NOR2_X1 U94 ( .A1(n14), .A2(n58), .ZN(B[20]) );
  AOI21_X1 U95 ( .B1(n114), .B2(n115), .A(SH[7]), .ZN(B[1]) );
  NAND2_X1 U96 ( .A1(n91), .A2(n116), .ZN(n115) );
  OAI221_X1 U97 ( .B1(n6), .B2(n55), .C1(n94), .C2(n56), .A(n117), .ZN(n116)
         );
  AOI22_X1 U98 ( .A1(A[2]), .A2(n1), .B1(A[1]), .B2(n7), .ZN(n117) );
  MUX2_X1 U99 ( .A(n118), .B(n119), .S(n86), .Z(n114) );
  AOI222_X1 U100 ( .A1(n100), .A2(n81), .B1(n101), .B2(n80), .C1(n103), .C2(
        n78), .ZN(n119) );
  OAI221_X1 U101 ( .B1(n5), .B2(n47), .C1(n4), .C2(n48), .A(n120), .ZN(n80) );
  AOI22_X1 U102 ( .A1(A[10]), .A2(n96), .B1(A[9]), .B2(n7), .ZN(n120) );
  OAI221_X1 U103 ( .B1(n93), .B2(n51), .C1(n3), .C2(n52), .A(n121), .ZN(n81)
         );
  AOI22_X1 U104 ( .A1(A[6]), .A2(n2), .B1(A[5]), .B2(n7), .ZN(n121) );
  NOR3_X1 U105 ( .A1(n12), .A2(n105), .A3(n122), .ZN(B[19]) );
  NOR2_X1 U106 ( .A1(n122), .A2(n110), .ZN(B[18]) );
  OR2_X1 U107 ( .A1(n12), .A2(n123), .ZN(n110) );
  NOR2_X1 U108 ( .A1(n122), .A2(n118), .ZN(B[17]) );
  OR2_X1 U109 ( .A1(n12), .A2(n59), .ZN(n118) );
  MUX2_X1 U110 ( .A(n79), .B(n29), .S(n13), .Z(n59) );
  NOR2_X1 U111 ( .A1(n122), .A2(n124), .ZN(B[16]) );
  OAI222_X1 U112 ( .A1(n23), .A2(n58), .B1(n69), .B2(n9), .C1(n26), .C2(n61), 
        .ZN(B[15]) );
  OAI222_X1 U113 ( .A1(n22), .A2(n58), .B1(n74), .B2(n9), .C1(n21), .C2(n61), 
        .ZN(B[14]) );
  OAI222_X1 U114 ( .A1(n27), .A2(n58), .B1(n79), .B2(n9), .C1(n29), .C2(n61), 
        .ZN(B[13]) );
  OAI221_X1 U115 ( .B1(n6), .B2(n39), .C1(n94), .C2(n40), .A(n125), .ZN(n77)
         );
  AOI22_X1 U116 ( .A1(A[18]), .A2(n1), .B1(A[17]), .B2(n7), .ZN(n125) );
  AOI222_X1 U117 ( .A1(n1), .A2(A[22]), .B1(n34), .B2(A[23]), .C1(n8), .C2(
        A[21]), .ZN(n79) );
  OAI221_X1 U118 ( .B1(n5), .B2(n43), .C1(n4), .C2(n44), .A(n126), .ZN(n78) );
  AOI22_X1 U119 ( .A1(A[14]), .A2(n96), .B1(A[13]), .B2(n7), .ZN(n126) );
  OAI222_X1 U120 ( .A1(n18), .A2(n58), .B1(n14), .B2(n9), .C1(n15), .C2(n61), 
        .ZN(B[12]) );
  NOR2_X1 U121 ( .A1(n60), .A2(SH[2]), .ZN(n64) );
  OAI222_X1 U122 ( .A1(n23), .A2(n61), .B1(n24), .B2(n58), .C1(n105), .C2(n60), 
        .ZN(B[11]) );
  MUX2_X1 U123 ( .A(n69), .B(n26), .S(n13), .Z(n105) );
  OAI221_X1 U124 ( .B1(n37), .B2(n93), .C1(n3), .C2(n38), .A(n127), .ZN(n67)
         );
  AOI22_X1 U125 ( .A1(A[20]), .A2(n2), .B1(A[19]), .B2(n7), .ZN(n127) );
  NAND2_X1 U126 ( .A1(n8), .A2(A[23]), .ZN(n69) );
  OAI221_X1 U127 ( .B1(n93), .B2(n45), .C1(n94), .C2(n46), .A(n128), .ZN(n102)
         );
  AOI22_X1 U128 ( .A1(A[12]), .A2(n1), .B1(A[11]), .B2(n8), .ZN(n128) );
  OAI221_X1 U129 ( .B1(n6), .B2(n41), .C1(n4), .C2(n42), .A(n129), .ZN(n65) );
  AOI22_X1 U130 ( .A1(A[16]), .A2(n96), .B1(A[15]), .B2(n8), .ZN(n129) );
  OAI222_X1 U131 ( .A1(n19), .A2(n58), .B1(n123), .B2(n60), .C1(n22), .C2(n61), 
        .ZN(B[10]) );
  OAI221_X1 U132 ( .B1(n5), .B2(n42), .C1(n3), .C2(n43), .A(n130), .ZN(n73) );
  AOI22_X1 U133 ( .A1(A[15]), .A2(n2), .B1(A[14]), .B2(n8), .ZN(n130) );
  NAND2_X1 U134 ( .A1(n10), .A2(n12), .ZN(n60) );
  NAND2_X1 U135 ( .A1(n86), .A2(n11), .ZN(n122) );
  MUX2_X1 U136 ( .A(n74), .B(n21), .S(n13), .Z(n123) );
  OAI221_X1 U137 ( .B1(n38), .B2(n6), .C1(n94), .C2(n39), .A(n131), .ZN(n72)
         );
  AOI22_X1 U138 ( .A1(A[19]), .A2(n1), .B1(A[18]), .B2(n8), .ZN(n131) );
  AOI22_X1 U139 ( .A1(A[22]), .A2(n7), .B1(A[23]), .B2(n2), .ZN(n74) );
  OAI221_X1 U140 ( .B1(n93), .B2(n46), .C1(n4), .C2(n47), .A(n132), .ZN(n112)
         );
  AOI22_X1 U141 ( .A1(A[11]), .A2(n96), .B1(A[10]), .B2(n8), .ZN(n132) );
  AOI21_X1 U142 ( .B1(n133), .B2(n134), .A(SH[7]), .ZN(B[0]) );
  NAND2_X1 U143 ( .A1(n91), .A2(n135), .ZN(n134) );
  OAI221_X1 U144 ( .B1(n6), .B2(n56), .C1(n3), .C2(n57), .A(n136), .ZN(n135)
         );
  AOI22_X1 U145 ( .A1(A[1]), .A2(n2), .B1(A[0]), .B2(n8), .ZN(n136) );
  AND3_X1 U146 ( .A1(n86), .A2(n13), .A3(n137), .ZN(n91) );
  MUX2_X1 U147 ( .A(n124), .B(n138), .S(n86), .Z(n133) );
  NOR2_X1 U148 ( .A1(SH[4]), .A2(n139), .ZN(n86) );
  AOI222_X1 U149 ( .A1(n100), .A2(n88), .B1(n101), .B2(n87), .C1(n103), .C2(
        n85), .ZN(n138) );
  OAI221_X1 U150 ( .B1(n5), .B2(n44), .C1(n94), .C2(n45), .A(n140), .ZN(n85)
         );
  AOI22_X1 U151 ( .A1(A[13]), .A2(n1), .B1(A[12]), .B2(n8), .ZN(n140) );
  NOR2_X1 U152 ( .A1(n13), .A2(n137), .ZN(n103) );
  OAI221_X1 U153 ( .B1(n93), .B2(n48), .C1(n4), .C2(n49), .A(n141), .ZN(n87)
         );
  AOI22_X1 U154 ( .A1(A[9]), .A2(n96), .B1(A[8]), .B2(n8), .ZN(n141) );
  NOR2_X1 U155 ( .A1(SH[2]), .A2(n137), .ZN(n101) );
  OAI221_X1 U156 ( .B1(n6), .B2(n52), .C1(n3), .C2(n53), .A(n142), .ZN(n88) );
  AOI22_X1 U157 ( .A1(A[5]), .A2(n2), .B1(A[4]), .B2(n8), .ZN(n142) );
  NOR2_X1 U158 ( .A1(n12), .A2(n13), .ZN(n100) );
  OR2_X1 U159 ( .A1(n12), .A2(n62), .ZN(n124) );
  MUX2_X1 U160 ( .A(n14), .B(n15), .S(n13), .Z(n62) );
  OAI221_X1 U161 ( .B1(n5), .B2(n40), .C1(n4), .C2(n41), .A(n143), .ZN(n84) );
  AOI22_X1 U162 ( .A1(A[17]), .A2(n1), .B1(A[16]), .B2(n8), .ZN(n143) );
  OAI221_X1 U163 ( .B1(n36), .B2(n5), .C1(n3), .C2(n37), .A(n144), .ZN(n83) );
  AOI22_X1 U164 ( .A1(A[21]), .A2(n96), .B1(A[20]), .B2(n7), .ZN(n144) );
  NOR2_X1 U165 ( .A1(SH[0]), .A2(SH[1]), .ZN(n97) );
  NOR2_X1 U166 ( .A1(n35), .A2(SH[1]), .ZN(n96) );
  NAND2_X1 U167 ( .A1(n35), .A2(SH[1]), .ZN(n94) );
  NAND2_X1 U168 ( .A1(SH[0]), .A2(SH[1]), .ZN(n93) );
  NOR2_X1 U169 ( .A1(SH[3]), .A2(n139), .ZN(n137) );
  OR2_X1 U170 ( .A1(SH[5]), .A2(SH[6]), .ZN(n139) );
endmodule


module fpAdder_DW01_sub_3 ( A, B, CI, DIFF, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9;
  wire   [7:1] carry;

  FA_X1 U2_7 ( .A(A[7]), .B(n2), .CI(carry[7]), .S(DIFF[7]) );
  FA_X1 U2_6 ( .A(A[6]), .B(n3), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  FA_X1 U2_5 ( .A(A[5]), .B(n4), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  FA_X1 U2_4 ( .A(A[4]), .B(n5), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  FA_X1 U2_3 ( .A(A[3]), .B(n6), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  FA_X1 U2_2 ( .A(A[2]), .B(n7), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  FA_X1 U2_1 ( .A(A[1]), .B(n8), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  INV_X1 U1 ( .A(B[7]), .ZN(n2) );
  XNOR2_X1 U2 ( .A(n9), .B(A[0]), .ZN(DIFF[0]) );
  INV_X1 U3 ( .A(B[1]), .ZN(n8) );
  NAND2_X1 U4 ( .A1(B[0]), .A2(n1), .ZN(carry[1]) );
  INV_X1 U5 ( .A(A[0]), .ZN(n1) );
  INV_X1 U6 ( .A(B[2]), .ZN(n7) );
  INV_X1 U7 ( .A(B[3]), .ZN(n6) );
  INV_X1 U8 ( .A(B[4]), .ZN(n5) );
  INV_X1 U9 ( .A(B[5]), .ZN(n4) );
  INV_X1 U10 ( .A(B[0]), .ZN(n9) );
  INV_X1 U11 ( .A(B[6]), .ZN(n3) );
endmodule


module fpAdder_DW_rash_1 ( A, DATA_TC, SH, SH_TC, B );
  input [23:0] A;
  input [7:0] SH;
  output [23:0] B;
  input DATA_TC, SH_TC;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144;

  NAND2_X1 U3 ( .A1(n100), .A2(n10), .ZN(n61) );
  INV_X1 U4 ( .A(n122), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n91), .A2(n11), .ZN(n58) );
  BUF_X1 U6 ( .A(n97), .Z(n7) );
  BUF_X1 U7 ( .A(n97), .Z(n8) );
  INV_X1 U8 ( .A(n137), .ZN(n12) );
  INV_X1 U9 ( .A(n64), .ZN(n9) );
  INV_X1 U10 ( .A(n69), .ZN(n25) );
  INV_X1 U11 ( .A(n79), .ZN(n28) );
  INV_X1 U12 ( .A(n74), .ZN(n20) );
  INV_X1 U13 ( .A(SH[2]), .ZN(n13) );
  INV_X1 U14 ( .A(SH[0]), .ZN(n35) );
  INV_X1 U15 ( .A(n83), .ZN(n14) );
  INV_X1 U16 ( .A(SH[7]), .ZN(n11) );
  INV_X1 U17 ( .A(n87), .ZN(n17) );
  INV_X1 U18 ( .A(n80), .ZN(n31) );
  INV_X1 U19 ( .A(n77), .ZN(n29) );
  INV_X1 U20 ( .A(n84), .ZN(n15) );
  INV_X1 U21 ( .A(n72), .ZN(n21) );
  INV_X1 U22 ( .A(n67), .ZN(n26) );
  INV_X1 U23 ( .A(n65), .ZN(n23) );
  INV_X1 U24 ( .A(n85), .ZN(n18) );
  INV_X1 U25 ( .A(n78), .ZN(n27) );
  INV_X1 U26 ( .A(n73), .ZN(n22) );
  INV_X1 U27 ( .A(n102), .ZN(n24) );
  INV_X1 U28 ( .A(n112), .ZN(n19) );
  INV_X1 U29 ( .A(n94), .ZN(n34) );
  INV_X1 U30 ( .A(n81), .ZN(n30) );
  INV_X1 U31 ( .A(n70), .ZN(n33) );
  INV_X1 U32 ( .A(n88), .ZN(n16) );
  INV_X1 U33 ( .A(n75), .ZN(n32) );
  INV_X1 U34 ( .A(A[23]), .ZN(n36) );
  INV_X1 U35 ( .A(A[2]), .ZN(n57) );
  INV_X1 U36 ( .A(A[22]), .ZN(n37) );
  INV_X1 U37 ( .A(A[21]), .ZN(n38) );
  INV_X1 U38 ( .A(A[19]), .ZN(n40) );
  INV_X1 U39 ( .A(A[20]), .ZN(n39) );
  INV_X1 U40 ( .A(A[11]), .ZN(n48) );
  INV_X1 U41 ( .A(A[12]), .ZN(n47) );
  INV_X1 U42 ( .A(A[18]), .ZN(n41) );
  INV_X1 U43 ( .A(A[3]), .ZN(n56) );
  INV_X1 U44 ( .A(A[14]), .ZN(n45) );
  INV_X1 U45 ( .A(A[10]), .ZN(n49) );
  INV_X1 U46 ( .A(A[6]), .ZN(n53) );
  INV_X1 U47 ( .A(A[15]), .ZN(n44) );
  INV_X1 U48 ( .A(A[7]), .ZN(n52) );
  INV_X1 U49 ( .A(A[16]), .ZN(n43) );
  INV_X1 U50 ( .A(A[8]), .ZN(n51) );
  INV_X1 U51 ( .A(A[17]), .ZN(n42) );
  INV_X1 U52 ( .A(A[4]), .ZN(n55) );
  INV_X1 U53 ( .A(A[13]), .ZN(n46) );
  INV_X1 U54 ( .A(A[5]), .ZN(n54) );
  INV_X1 U55 ( .A(A[9]), .ZN(n50) );
  NOR2_X1 U56 ( .A1(n35), .A2(SH[1]), .ZN(n1) );
  NOR2_X1 U57 ( .A1(n35), .A2(SH[1]), .ZN(n2) );
  NAND2_X1 U58 ( .A1(n35), .A2(SH[1]), .ZN(n3) );
  NAND2_X1 U59 ( .A1(n35), .A2(SH[1]), .ZN(n4) );
  NAND2_X1 U60 ( .A1(SH[0]), .A2(SH[1]), .ZN(n5) );
  NAND2_X1 U61 ( .A1(SH[0]), .A2(SH[1]), .ZN(n6) );
  OAI222_X1 U62 ( .A1(n31), .A2(n58), .B1(n59), .B2(n60), .C1(n27), .C2(n61), 
        .ZN(B[9]) );
  OAI222_X1 U63 ( .A1(n17), .A2(n58), .B1(n62), .B2(n60), .C1(n18), .C2(n61), 
        .ZN(B[8]) );
  OAI221_X1 U64 ( .B1(n33), .B2(n58), .C1(n24), .C2(n61), .A(n63), .ZN(B[7])
         );
  AOI222_X1 U65 ( .A1(n64), .A2(n65), .B1(n66), .B2(n67), .C1(n68), .C2(n25), 
        .ZN(n63) );
  OAI221_X1 U66 ( .B1(n32), .B2(n58), .C1(n19), .C2(n61), .A(n71), .ZN(B[6])
         );
  AOI222_X1 U67 ( .A1(n68), .A2(n20), .B1(n66), .B2(n72), .C1(n64), .C2(n73), 
        .ZN(n71) );
  OAI221_X1 U68 ( .B1(n30), .B2(n58), .C1(n31), .C2(n61), .A(n76), .ZN(B[5])
         );
  AOI222_X1 U69 ( .A1(n68), .A2(n28), .B1(n66), .B2(n77), .C1(n64), .C2(n78), 
        .ZN(n76) );
  OAI221_X1 U70 ( .B1(n16), .B2(n58), .C1(n17), .C2(n61), .A(n82), .ZN(B[4])
         );
  AOI222_X1 U71 ( .A1(n68), .A2(n83), .B1(n66), .B2(n84), .C1(n64), .C2(n85), 
        .ZN(n82) );
  NOR2_X1 U72 ( .A1(n60), .A2(n13), .ZN(n66) );
  NOR4_X1 U73 ( .A1(n12), .A2(SH[2]), .A3(n86), .A4(SH[7]), .ZN(n68) );
  AOI21_X1 U74 ( .B1(n89), .B2(n90), .A(SH[7]), .ZN(B[3]) );
  NAND2_X1 U75 ( .A1(n91), .A2(n92), .ZN(n90) );
  OAI221_X1 U76 ( .B1(n93), .B2(n53), .C1(n3), .C2(n54), .A(n95), .ZN(n92) );
  AOI22_X1 U77 ( .A1(A[4]), .A2(n2), .B1(A[3]), .B2(n7), .ZN(n95) );
  MUX2_X1 U78 ( .A(n98), .B(n99), .S(n86), .Z(n89) );
  AOI222_X1 U79 ( .A1(n100), .A2(n70), .B1(n101), .B2(n102), .C1(n103), .C2(
        n65), .ZN(n99) );
  OAI221_X1 U80 ( .B1(n6), .B2(n49), .C1(n94), .C2(n50), .A(n104), .ZN(n70) );
  AOI22_X1 U81 ( .A1(A[8]), .A2(n1), .B1(A[7]), .B2(n7), .ZN(n104) );
  OR2_X1 U82 ( .A1(n12), .A2(n105), .ZN(n98) );
  AOI21_X1 U83 ( .B1(n106), .B2(n107), .A(SH[7]), .ZN(B[2]) );
  NAND2_X1 U84 ( .A1(n91), .A2(n108), .ZN(n107) );
  OAI221_X1 U85 ( .B1(n5), .B2(n54), .C1(n4), .C2(n55), .A(n109), .ZN(n108) );
  AOI22_X1 U86 ( .A1(A[3]), .A2(n96), .B1(A[2]), .B2(n7), .ZN(n109) );
  MUX2_X1 U87 ( .A(n110), .B(n111), .S(n86), .Z(n106) );
  AOI222_X1 U88 ( .A1(n100), .A2(n75), .B1(n101), .B2(n112), .C1(n103), .C2(
        n73), .ZN(n111) );
  OAI221_X1 U89 ( .B1(n93), .B2(n50), .C1(n3), .C2(n51), .A(n113), .ZN(n75) );
  AOI22_X1 U90 ( .A1(A[7]), .A2(n2), .B1(A[6]), .B2(n7), .ZN(n113) );
  NOR2_X1 U91 ( .A1(n58), .A2(n69), .ZN(B[23]) );
  NOR2_X1 U92 ( .A1(n74), .A2(n58), .ZN(B[22]) );
  NOR2_X1 U93 ( .A1(n79), .A2(n58), .ZN(B[21]) );
  NOR2_X1 U94 ( .A1(n14), .A2(n58), .ZN(B[20]) );
  AOI21_X1 U95 ( .B1(n114), .B2(n115), .A(SH[7]), .ZN(B[1]) );
  NAND2_X1 U96 ( .A1(n91), .A2(n116), .ZN(n115) );
  OAI221_X1 U97 ( .B1(n6), .B2(n55), .C1(n94), .C2(n56), .A(n117), .ZN(n116)
         );
  AOI22_X1 U98 ( .A1(A[2]), .A2(n1), .B1(A[1]), .B2(n7), .ZN(n117) );
  MUX2_X1 U99 ( .A(n118), .B(n119), .S(n86), .Z(n114) );
  AOI222_X1 U100 ( .A1(n100), .A2(n81), .B1(n101), .B2(n80), .C1(n103), .C2(
        n78), .ZN(n119) );
  OAI221_X1 U101 ( .B1(n5), .B2(n47), .C1(n4), .C2(n48), .A(n120), .ZN(n80) );
  AOI22_X1 U102 ( .A1(A[10]), .A2(n96), .B1(A[9]), .B2(n7), .ZN(n120) );
  OAI221_X1 U103 ( .B1(n93), .B2(n51), .C1(n3), .C2(n52), .A(n121), .ZN(n81)
         );
  AOI22_X1 U104 ( .A1(A[6]), .A2(n2), .B1(A[5]), .B2(n7), .ZN(n121) );
  NOR3_X1 U105 ( .A1(n12), .A2(n105), .A3(n122), .ZN(B[19]) );
  NOR2_X1 U106 ( .A1(n122), .A2(n110), .ZN(B[18]) );
  OR2_X1 U107 ( .A1(n12), .A2(n123), .ZN(n110) );
  NOR2_X1 U108 ( .A1(n122), .A2(n118), .ZN(B[17]) );
  OR2_X1 U109 ( .A1(n12), .A2(n59), .ZN(n118) );
  MUX2_X1 U110 ( .A(n79), .B(n29), .S(n13), .Z(n59) );
  NOR2_X1 U111 ( .A1(n122), .A2(n124), .ZN(B[16]) );
  OAI222_X1 U112 ( .A1(n23), .A2(n58), .B1(n69), .B2(n9), .C1(n26), .C2(n61), 
        .ZN(B[15]) );
  OAI222_X1 U113 ( .A1(n22), .A2(n58), .B1(n74), .B2(n9), .C1(n21), .C2(n61), 
        .ZN(B[14]) );
  OAI222_X1 U114 ( .A1(n27), .A2(n58), .B1(n79), .B2(n9), .C1(n29), .C2(n61), 
        .ZN(B[13]) );
  OAI221_X1 U115 ( .B1(n6), .B2(n39), .C1(n94), .C2(n40), .A(n125), .ZN(n77)
         );
  AOI22_X1 U116 ( .A1(A[18]), .A2(n1), .B1(A[17]), .B2(n7), .ZN(n125) );
  AOI222_X1 U117 ( .A1(n1), .A2(A[22]), .B1(n34), .B2(A[23]), .C1(n8), .C2(
        A[21]), .ZN(n79) );
  OAI221_X1 U118 ( .B1(n5), .B2(n43), .C1(n4), .C2(n44), .A(n126), .ZN(n78) );
  AOI22_X1 U119 ( .A1(A[14]), .A2(n96), .B1(A[13]), .B2(n7), .ZN(n126) );
  OAI222_X1 U120 ( .A1(n18), .A2(n58), .B1(n14), .B2(n9), .C1(n15), .C2(n61), 
        .ZN(B[12]) );
  NOR2_X1 U121 ( .A1(n60), .A2(SH[2]), .ZN(n64) );
  OAI222_X1 U122 ( .A1(n23), .A2(n61), .B1(n24), .B2(n58), .C1(n105), .C2(n60), 
        .ZN(B[11]) );
  MUX2_X1 U123 ( .A(n69), .B(n26), .S(n13), .Z(n105) );
  OAI221_X1 U124 ( .B1(n37), .B2(n93), .C1(n3), .C2(n38), .A(n127), .ZN(n67)
         );
  AOI22_X1 U125 ( .A1(A[20]), .A2(n2), .B1(A[19]), .B2(n7), .ZN(n127) );
  NAND2_X1 U126 ( .A1(n8), .A2(A[23]), .ZN(n69) );
  OAI221_X1 U127 ( .B1(n93), .B2(n45), .C1(n94), .C2(n46), .A(n128), .ZN(n102)
         );
  AOI22_X1 U128 ( .A1(A[12]), .A2(n1), .B1(A[11]), .B2(n8), .ZN(n128) );
  OAI221_X1 U129 ( .B1(n6), .B2(n41), .C1(n4), .C2(n42), .A(n129), .ZN(n65) );
  AOI22_X1 U130 ( .A1(A[16]), .A2(n96), .B1(A[15]), .B2(n8), .ZN(n129) );
  OAI222_X1 U131 ( .A1(n19), .A2(n58), .B1(n123), .B2(n60), .C1(n22), .C2(n61), 
        .ZN(B[10]) );
  OAI221_X1 U132 ( .B1(n5), .B2(n42), .C1(n3), .C2(n43), .A(n130), .ZN(n73) );
  AOI22_X1 U133 ( .A1(A[15]), .A2(n2), .B1(A[14]), .B2(n8), .ZN(n130) );
  NAND2_X1 U134 ( .A1(n10), .A2(n12), .ZN(n60) );
  NAND2_X1 U135 ( .A1(n86), .A2(n11), .ZN(n122) );
  MUX2_X1 U136 ( .A(n74), .B(n21), .S(n13), .Z(n123) );
  OAI221_X1 U137 ( .B1(n38), .B2(n6), .C1(n94), .C2(n39), .A(n131), .ZN(n72)
         );
  AOI22_X1 U138 ( .A1(A[19]), .A2(n1), .B1(A[18]), .B2(n8), .ZN(n131) );
  AOI22_X1 U139 ( .A1(A[22]), .A2(n7), .B1(A[23]), .B2(n2), .ZN(n74) );
  OAI221_X1 U140 ( .B1(n93), .B2(n46), .C1(n4), .C2(n47), .A(n132), .ZN(n112)
         );
  AOI22_X1 U141 ( .A1(A[11]), .A2(n96), .B1(A[10]), .B2(n8), .ZN(n132) );
  AOI21_X1 U142 ( .B1(n133), .B2(n134), .A(SH[7]), .ZN(B[0]) );
  NAND2_X1 U143 ( .A1(n91), .A2(n135), .ZN(n134) );
  OAI221_X1 U144 ( .B1(n6), .B2(n56), .C1(n3), .C2(n57), .A(n136), .ZN(n135)
         );
  AOI22_X1 U145 ( .A1(A[1]), .A2(n2), .B1(A[0]), .B2(n8), .ZN(n136) );
  AND3_X1 U146 ( .A1(n86), .A2(n13), .A3(n137), .ZN(n91) );
  MUX2_X1 U147 ( .A(n124), .B(n138), .S(n86), .Z(n133) );
  NOR2_X1 U148 ( .A1(SH[4]), .A2(n139), .ZN(n86) );
  AOI222_X1 U149 ( .A1(n100), .A2(n88), .B1(n101), .B2(n87), .C1(n103), .C2(
        n85), .ZN(n138) );
  OAI221_X1 U150 ( .B1(n5), .B2(n44), .C1(n94), .C2(n45), .A(n140), .ZN(n85)
         );
  AOI22_X1 U151 ( .A1(A[13]), .A2(n1), .B1(A[12]), .B2(n8), .ZN(n140) );
  NOR2_X1 U152 ( .A1(n13), .A2(n137), .ZN(n103) );
  OAI221_X1 U153 ( .B1(n93), .B2(n48), .C1(n4), .C2(n49), .A(n141), .ZN(n87)
         );
  AOI22_X1 U154 ( .A1(A[9]), .A2(n96), .B1(A[8]), .B2(n8), .ZN(n141) );
  NOR2_X1 U155 ( .A1(SH[2]), .A2(n137), .ZN(n101) );
  OAI221_X1 U156 ( .B1(n6), .B2(n52), .C1(n3), .C2(n53), .A(n142), .ZN(n88) );
  AOI22_X1 U157 ( .A1(A[5]), .A2(n2), .B1(A[4]), .B2(n8), .ZN(n142) );
  NOR2_X1 U158 ( .A1(n12), .A2(n13), .ZN(n100) );
  OR2_X1 U159 ( .A1(n12), .A2(n62), .ZN(n124) );
  MUX2_X1 U160 ( .A(n14), .B(n15), .S(n13), .Z(n62) );
  OAI221_X1 U161 ( .B1(n5), .B2(n40), .C1(n4), .C2(n41), .A(n143), .ZN(n84) );
  AOI22_X1 U162 ( .A1(A[17]), .A2(n1), .B1(A[16]), .B2(n8), .ZN(n143) );
  OAI221_X1 U163 ( .B1(n36), .B2(n5), .C1(n3), .C2(n37), .A(n144), .ZN(n83) );
  AOI22_X1 U164 ( .A1(A[21]), .A2(n96), .B1(A[20]), .B2(n7), .ZN(n144) );
  NOR2_X1 U165 ( .A1(SH[0]), .A2(SH[1]), .ZN(n97) );
  NOR2_X1 U166 ( .A1(n35), .A2(SH[1]), .ZN(n96) );
  NAND2_X1 U167 ( .A1(n35), .A2(SH[1]), .ZN(n94) );
  NAND2_X1 U168 ( .A1(SH[0]), .A2(SH[1]), .ZN(n93) );
  NOR2_X1 U169 ( .A1(SH[3]), .A2(n139), .ZN(n137) );
  OR2_X1 U170 ( .A1(SH[5]), .A2(SH[6]), .ZN(n139) );
endmodule


module fpAdder_DW01_sub_4 ( A, B, CI, DIFF, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9;
  wire   [7:1] carry;

  FA_X1 U2_7 ( .A(A[7]), .B(n2), .CI(carry[7]), .S(DIFF[7]) );
  FA_X1 U2_6 ( .A(A[6]), .B(n3), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  FA_X1 U2_5 ( .A(A[5]), .B(n4), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  FA_X1 U2_4 ( .A(A[4]), .B(n5), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  FA_X1 U2_3 ( .A(A[3]), .B(n6), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  FA_X1 U2_2 ( .A(A[2]), .B(n7), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  FA_X1 U2_1 ( .A(A[1]), .B(n8), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  INV_X1 U1 ( .A(B[7]), .ZN(n2) );
  XNOR2_X1 U2 ( .A(n9), .B(A[0]), .ZN(DIFF[0]) );
  INV_X1 U3 ( .A(B[1]), .ZN(n8) );
  NAND2_X1 U4 ( .A1(B[0]), .A2(n1), .ZN(carry[1]) );
  INV_X1 U5 ( .A(A[0]), .ZN(n1) );
  INV_X1 U6 ( .A(B[2]), .ZN(n7) );
  INV_X1 U7 ( .A(B[3]), .ZN(n6) );
  INV_X1 U8 ( .A(B[4]), .ZN(n5) );
  INV_X1 U9 ( .A(B[5]), .ZN(n4) );
  INV_X1 U10 ( .A(B[0]), .ZN(n9) );
  INV_X1 U11 ( .A(B[6]), .ZN(n3) );
endmodule


module fpAdder_DW01_sub_5 ( A, B, CI, DIFF, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7;
  wire   [7:1] carry;

  FA_X1 U2_7 ( .A(A[7]), .B(n2), .CI(carry[7]), .S(DIFF[7]) );
  FA_X1 U2_6 ( .A(A[6]), .B(n2), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  FA_X1 U2_5 ( .A(A[5]), .B(n2), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  FA_X1 U2_4 ( .A(A[4]), .B(n3), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  FA_X1 U2_3 ( .A(A[3]), .B(n4), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  FA_X1 U2_2 ( .A(A[2]), .B(n5), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  FA_X1 U2_1 ( .A(A[1]), .B(n6), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  INV_X1 U1 ( .A(B[5]), .ZN(n2) );
  XNOR2_X1 U2 ( .A(n7), .B(A[0]), .ZN(DIFF[0]) );
  INV_X1 U3 ( .A(B[4]), .ZN(n3) );
  INV_X1 U4 ( .A(B[3]), .ZN(n4) );
  INV_X1 U5 ( .A(B[2]), .ZN(n5) );
  INV_X1 U6 ( .A(B[1]), .ZN(n6) );
  NAND2_X1 U7 ( .A1(B[0]), .A2(n1), .ZN(carry[1]) );
  INV_X1 U8 ( .A(B[0]), .ZN(n7) );
  INV_X1 U9 ( .A(A[0]), .ZN(n1) );
endmodule


module fpAdder ( clk, reset, enable, A, B, result, overFlow );
  input [31:0] A;
  input [31:0] B;
  output [31:0] result;
  input clk, reset, enable;
  output overFlow;
  wire   IBA, IBB, N135, N137, N138, N139, N140, N141, N142, N143, N144, N145,
         N146, N147, N148, N149, N150, N151, N152, N153, N154, N155, N156,
         N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167,
         N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178,
         N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189,
         N190, N191, N192, N193, N194, N195, N196, N197, N198, N199, N200,
         N201, N202, N203, N204, N205, N206, N207, N208, N212, N213, N214,
         N215, N216, N217, N218, N219, N220, N221, N222, N223, N224, N225,
         N226, N227, N228, N229, N230, N231, N232, N233, N234, N235, N236,
         N238, N239, N240, N241, N242, N243, N244, N245, N278, N280, N281,
         N282, N283, N284, N285, N286, N287, N288, N289, N290, N291, N292,
         N293, N294, N295, N296, N297, N298, N299, N300, N301, N302, N303,
         N304, N305, N306, N307, N308, N309, N310, N311, N312, N313, N314,
         N315, N316, N317, N318, N319, N320, N321, N322, N323, N324, N325,
         N326, N327, N480, N481, N482, N483, N484, N517, N518, N521, N549,
         N550, N551, N552, N553, N554, N555, N556, N557, N558, N559, N560,
         N561, N562, N563, N564, N565, N566, N567, N568, N569, N570, N571,
         N580, N581, N582, N583, N584, N585, N586, N587, N612, n74, n1350,
         n1410, n1420, n1430, n1440, n1450, n1460, n1470, n1480, n1490, n1500,
         n1510, n1520, n1530, n1540, n1550, n1560, n1570, n1580, n1590, n1600,
         n1610, n1620, n1630, n1640, n1650, n1720, n1730, n1740, n1750, n1760,
         n1770, n1780, n1790, n1800, n1810, n1820, n1830, n1840, n1850, n1860,
         n1870, n1880, n1890, n1900, n1910, n1920, n1930, n1940, n1950, n1960,
         n1980, n1990, n2000, n2010, n2020, n2030, n2040, n2050, n2060, n2070,
         n2080, n209, n210, n211, n2120, n2130, n2140, n2150, n2160, n2170,
         n2180, n2190, n2200, n2210, n2220, n2230, n2240, n2250, n2260, n2270,
         n2280, n2290, n2300, n2310, n2320, n2330, n2340, n2350, n2360, n237,
         n2380, n2390, n2400, n2410, n2420, n2430, n2440, n2450, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n2780, n279, n2800,
         n2810, n2820, n2830, n2840, n2850, n2860, n2870, n2880, n2890, n2900,
         n2910, n2920, n2930, n2940, n2950, n2960, n2970, n2980, n2990, n3000,
         n3010, n3020, n3030, n3040, n3050, n3060, n3070, n3080, n3090, n3100,
         n3110, n3120, n3130, n3140, n3150, n3160, n3170, n3180, n3190, n3200,
         n3210, n3220, n3230, n3240, n3250, n3260, n3270, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n4800, n4810, n4820, n4830, n4840,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, N576,
         N575, N574, r145_B_23_, sll_78_ML_int_5__16_, sll_78_ML_int_5__17_,
         sll_78_ML_int_5__18_, sll_78_ML_int_5__19_, sll_78_ML_int_5__20_,
         sll_78_ML_int_5__21_, sll_78_ML_int_5__22_, sll_78_ML_int_4__8_,
         sll_78_ML_int_4__9_, sll_78_ML_int_4__10_, sll_78_ML_int_4__11_,
         sll_78_ML_int_4__12_, sll_78_ML_int_4__13_, sll_78_ML_int_4__14_,
         sll_78_ML_int_4__15_, sll_78_ML_int_4__16_, sll_78_ML_int_4__17_,
         sll_78_ML_int_4__18_, sll_78_ML_int_4__19_, sll_78_ML_int_4__20_,
         sll_78_ML_int_4__21_, sll_78_ML_int_4__22_, sll_78_ML_int_3__0_,
         sll_78_ML_int_3__1_, sll_78_ML_int_3__2_, sll_78_ML_int_3__3_,
         sll_78_ML_int_3__4_, sll_78_ML_int_3__5_, sll_78_ML_int_3__6_,
         sll_78_ML_int_3__7_, sll_78_ML_int_3__8_, sll_78_ML_int_3__9_,
         sll_78_ML_int_3__10_, sll_78_ML_int_3__11_, sll_78_ML_int_3__12_,
         sll_78_ML_int_3__13_, sll_78_ML_int_3__14_, sll_78_ML_int_3__15_,
         sll_78_ML_int_3__16_, sll_78_ML_int_3__17_, sll_78_ML_int_3__18_,
         sll_78_ML_int_3__19_, sll_78_ML_int_3__20_, sll_78_ML_int_3__21_,
         sll_78_ML_int_3__22_, sll_78_ML_int_2__0_, sll_78_ML_int_2__1_,
         sll_78_ML_int_2__2_, sll_78_ML_int_2__3_, sll_78_ML_int_2__4_,
         sll_78_ML_int_2__5_, sll_78_ML_int_2__6_, sll_78_ML_int_2__7_,
         sll_78_ML_int_2__8_, sll_78_ML_int_2__9_, sll_78_ML_int_2__10_,
         sll_78_ML_int_2__11_, sll_78_ML_int_2__12_, sll_78_ML_int_2__13_,
         sll_78_ML_int_2__14_, sll_78_ML_int_2__15_, sll_78_ML_int_2__16_,
         sll_78_ML_int_2__17_, sll_78_ML_int_2__18_, sll_78_ML_int_2__19_,
         sll_78_ML_int_2__20_, sll_78_ML_int_2__21_, sll_78_ML_int_2__22_,
         sll_78_ML_int_1__0_, sll_78_ML_int_1__1_, sll_78_ML_int_1__2_,
         sll_78_ML_int_1__3_, sll_78_ML_int_1__4_, sll_78_ML_int_1__5_,
         sll_78_ML_int_1__6_, sll_78_ML_int_1__7_, sll_78_ML_int_1__8_,
         sll_78_ML_int_1__9_, sll_78_ML_int_1__10_, sll_78_ML_int_1__11_,
         sll_78_ML_int_1__12_, sll_78_ML_int_1__13_, sll_78_ML_int_1__14_,
         sll_78_ML_int_1__15_, sll_78_ML_int_1__16_, sll_78_ML_int_1__17_,
         sll_78_ML_int_1__18_, sll_78_ML_int_1__19_, sll_78_ML_int_1__20_,
         sll_78_ML_int_1__21_, sll_78_ML_int_1__22_, sll_78_A_0_, sll_78_A_1_,
         sll_78_A_2_, sll_78_A_3_, sll_78_A_4_, sll_78_A_5_, sll_78_A_6_,
         sll_78_A_7_, sll_78_A_8_, sll_78_A_9_, sll_78_A_10_, sll_78_A_11_,
         sll_78_A_12_, sll_78_A_13_, sll_78_A_14_, sll_78_A_15_, sll_78_A_16_,
         sll_78_A_17_, sll_78_A_18_, sll_78_A_19_, sll_78_A_20_, sll_78_A_21_,
         sll_78_A_22_, sub_78_carry_5_, sub_78_B_0_, sub_78_B_1_, sub_78_B_2_,
         sub_78_B_4_, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n5170, n5180, n519, n520, n5210, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n5490, n5500, n5510, n5520, n5530, n5540, n5550, n5560, n5570,
         n5580, n5590, n5600, n5610, n5620, n5630, n5640, n5650, n5660, n5670,
         n5680, n5690, n5700, n5710, n572, n573, n5740, n5750, n5760, n577,
         n578, n579, n5800, n5810, n5820, n5830, n5840, n5850, n5860, n5870,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n6120, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749;
  wire   [30:0] A_reg;
  wire   [31:0] B_reg;
  wire   [23:0] MB;
  wire   [22:0] MA;
  wire   [4:0] MSB;

  DFF_X1 A_reg_reg_31_ ( .D(n473), .CK(clk), .QN(n1650) );
  DFF_X1 result_reg_31_ ( .D(n720), .CK(clk), .Q(result[31]) );
  DFF_X1 result_reg_30_ ( .D(n432), .CK(clk), .Q(result[30]) );
  DFF_X1 result_reg_29_ ( .D(n433), .CK(clk), .Q(result[29]) );
  DFF_X1 result_reg_28_ ( .D(n434), .CK(clk), .Q(result[28]) );
  DFF_X1 result_reg_27_ ( .D(n435), .CK(clk), .Q(result[27]) );
  DFF_X1 result_reg_26_ ( .D(n436), .CK(clk), .Q(result[26]) );
  DFF_X1 result_reg_25_ ( .D(n437), .CK(clk), .Q(result[25]) );
  DFF_X1 result_reg_24_ ( .D(n438), .CK(clk), .Q(result[24]) );
  DFF_X1 result_reg_23_ ( .D(n439), .CK(clk), .Q(result[23]) );
  DFF_X1 overFlow_reg ( .D(n441), .CK(clk), .Q(overFlow) );
  DLH_X1 MSB_reg_4_ ( .G(N612), .D(N484), .Q(MSB[4]) );
  DLH_X1 MSB_reg_3_ ( .G(N612), .D(N483), .Q(MSB[3]) );
  DLH_X1 MSB_reg_2_ ( .G(N612), .D(N482), .Q(MSB[2]) );
  DLH_X1 MSB_reg_1_ ( .G(N612), .D(N481), .Q(MSB[1]) );
  DLH_X1 MSB_reg_0_ ( .G(N612), .D(N480), .Q(MSB[0]) );
  DFF_X1 result_reg_0_ ( .D(n440), .CK(clk), .Q(result[0]) );
  DFF_X1 result_reg_1_ ( .D(n676), .CK(clk), .Q(result[1]) );
  DFF_X1 result_reg_2_ ( .D(n678), .CK(clk), .Q(result[2]) );
  DFF_X1 result_reg_3_ ( .D(n680), .CK(clk), .Q(result[3]) );
  DFF_X1 result_reg_4_ ( .D(n682), .CK(clk), .Q(result[4]) );
  DFF_X1 result_reg_5_ ( .D(n684), .CK(clk), .Q(result[5]) );
  DFF_X1 result_reg_6_ ( .D(n686), .CK(clk), .Q(result[6]) );
  DFF_X1 result_reg_7_ ( .D(n688), .CK(clk), .Q(result[7]) );
  DFF_X1 result_reg_8_ ( .D(n690), .CK(clk), .Q(result[8]) );
  DFF_X1 result_reg_9_ ( .D(n692), .CK(clk), .Q(result[9]) );
  DFF_X1 result_reg_10_ ( .D(n694), .CK(clk), .Q(result[10]) );
  DFF_X1 result_reg_11_ ( .D(n696), .CK(clk), .Q(result[11]) );
  DFF_X1 result_reg_12_ ( .D(n698), .CK(clk), .Q(result[12]) );
  DFF_X1 result_reg_13_ ( .D(n700), .CK(clk), .Q(result[13]) );
  DFF_X1 result_reg_14_ ( .D(n702), .CK(clk), .Q(result[14]) );
  DFF_X1 result_reg_15_ ( .D(n704), .CK(clk), .Q(result[15]) );
  DFF_X1 result_reg_16_ ( .D(n706), .CK(clk), .Q(result[16]) );
  DFF_X1 result_reg_17_ ( .D(n708), .CK(clk), .Q(result[17]) );
  DFF_X1 result_reg_18_ ( .D(n710), .CK(clk), .Q(result[18]) );
  DFF_X1 result_reg_19_ ( .D(n712), .CK(clk), .Q(result[19]) );
  DFF_X1 result_reg_20_ ( .D(n714), .CK(clk), .Q(result[20]) );
  DFF_X1 result_reg_21_ ( .D(n716), .CK(clk), .Q(result[21]) );
  DFF_X1 result_reg_22_ ( .D(n718), .CK(clk), .Q(result[22]) );
  fpAdder_DW01_sub_1 sub_70 ( .A(MB), .B({r145_B_23_, MA}), .CI(1'b0), .DIFF({
        N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, 
        N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304}) );
  fpAdder_DW01_sub_2 sub_68 ( .A({r145_B_23_, MA}), .B(MB), .CI(1'b0), .DIFF({
        N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, 
        N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280}) );
  fpAdder_DW01_inc_0 add_63 ( .A({N208, N207, N206, N205, N204, N203, N202, 
        N201}), .SUM({N245, N244, N243, N242, N241, N240, N239, N238}) );
  fpAdder_DW01_add_0 add_59 ( .A({1'b0, r145_B_23_, MA}), .B({1'b0, MB}), .CI(
        1'b0), .SUM({N236, N235, N234, N233, N232, N231, N230, N229, N228, 
        N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, 
        N215, N214, N213, N212}) );
  fpAdder_DW_rash_0 srl_52 ( .A({IBB, B_reg[22:0]}), .DATA_TC(1'b0), .SH({N144, 
        N143, N142, N141, N140, N139, N138, N137}), .SH_TC(1'b0), .B({N168, 
        N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, 
        N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145}) );
  fpAdder_DW01_sub_3 sub_52 ( .A(A_reg[30:23]), .B(B_reg[30:23]), .CI(1'b0), 
        .DIFF({N144, N143, N142, N141, N140, N139, N138, N137}) );
  fpAdder_DW_rash_1 srl_55 ( .A({IBA, A_reg[22:0]}), .DATA_TC(1'b0), .SH({N176, 
        N175, N174, N173, N172, N171, N170, N169}), .SH_TC(1'b0), .B({N200, 
        N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, 
        N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177}) );
  fpAdder_DW01_sub_4 sub_55 ( .A(B_reg[30:23]), .B(A_reg[30:23]), .CI(1'b0), 
        .DIFF({N176, N175, N174, N173, N172, N171, N170, N169}) );
  fpAdder_DW01_sub_5 sub_79_2 ( .A({N208, N207, N206, N205, N204, N203, N202, 
        N201}), .B({n506, n506, n506, N576, N575, N574, n344, n343}), .CI(1'b0), .DIFF({N587, N586, N585, N584, N583, N582, N581, N580}) );
  MUX2_X1 sll_78_M1_0_1 ( .A(sll_78_A_1_), .B(sll_78_A_0_), .S(N517), .Z(
        sll_78_ML_int_1__1_) );
  MUX2_X1 sll_78_M1_0_2 ( .A(sll_78_A_2_), .B(sll_78_A_1_), .S(N517), .Z(
        sll_78_ML_int_1__2_) );
  MUX2_X1 sll_78_M1_0_3 ( .A(sll_78_A_3_), .B(sll_78_A_2_), .S(N517), .Z(
        sll_78_ML_int_1__3_) );
  MUX2_X1 sll_78_M1_0_4 ( .A(sll_78_A_4_), .B(sll_78_A_3_), .S(N517), .Z(
        sll_78_ML_int_1__4_) );
  MUX2_X1 sll_78_M1_0_5 ( .A(sll_78_A_5_), .B(sll_78_A_4_), .S(N517), .Z(
        sll_78_ML_int_1__5_) );
  MUX2_X1 sll_78_M1_0_6 ( .A(sll_78_A_6_), .B(sll_78_A_5_), .S(N517), .Z(
        sll_78_ML_int_1__6_) );
  MUX2_X1 sll_78_M1_0_7 ( .A(sll_78_A_7_), .B(sll_78_A_6_), .S(N517), .Z(
        sll_78_ML_int_1__7_) );
  MUX2_X1 sll_78_M1_0_8 ( .A(sll_78_A_8_), .B(sll_78_A_7_), .S(N517), .Z(
        sll_78_ML_int_1__8_) );
  MUX2_X1 sll_78_M1_0_9 ( .A(sll_78_A_9_), .B(sll_78_A_8_), .S(N517), .Z(
        sll_78_ML_int_1__9_) );
  MUX2_X1 sll_78_M1_0_10 ( .A(sll_78_A_10_), .B(sll_78_A_9_), .S(N517), .Z(
        sll_78_ML_int_1__10_) );
  MUX2_X1 sll_78_M1_0_11 ( .A(sll_78_A_11_), .B(sll_78_A_10_), .S(N517), .Z(
        sll_78_ML_int_1__11_) );
  MUX2_X1 sll_78_M1_0_12 ( .A(sll_78_A_12_), .B(sll_78_A_11_), .S(N517), .Z(
        sll_78_ML_int_1__12_) );
  MUX2_X1 sll_78_M1_0_13 ( .A(sll_78_A_13_), .B(sll_78_A_12_), .S(N517), .Z(
        sll_78_ML_int_1__13_) );
  MUX2_X1 sll_78_M1_0_14 ( .A(sll_78_A_14_), .B(sll_78_A_13_), .S(N517), .Z(
        sll_78_ML_int_1__14_) );
  MUX2_X1 sll_78_M1_0_15 ( .A(sll_78_A_15_), .B(sll_78_A_14_), .S(N517), .Z(
        sll_78_ML_int_1__15_) );
  MUX2_X1 sll_78_M1_0_16 ( .A(sll_78_A_16_), .B(sll_78_A_15_), .S(N517), .Z(
        sll_78_ML_int_1__16_) );
  MUX2_X1 sll_78_M1_0_17 ( .A(sll_78_A_17_), .B(sll_78_A_16_), .S(N517), .Z(
        sll_78_ML_int_1__17_) );
  MUX2_X1 sll_78_M1_0_18 ( .A(sll_78_A_18_), .B(sll_78_A_17_), .S(N517), .Z(
        sll_78_ML_int_1__18_) );
  MUX2_X1 sll_78_M1_0_19 ( .A(sll_78_A_19_), .B(sll_78_A_18_), .S(N517), .Z(
        sll_78_ML_int_1__19_) );
  MUX2_X1 sll_78_M1_0_20 ( .A(sll_78_A_20_), .B(sll_78_A_19_), .S(N517), .Z(
        sll_78_ML_int_1__20_) );
  MUX2_X1 sll_78_M1_0_21 ( .A(sll_78_A_21_), .B(sll_78_A_20_), .S(N517), .Z(
        sll_78_ML_int_1__21_) );
  MUX2_X1 sll_78_M1_0_22 ( .A(sll_78_A_22_), .B(sll_78_A_21_), .S(N517), .Z(
        sll_78_ML_int_1__22_) );
  MUX2_X1 sll_78_M1_1_2 ( .A(sll_78_ML_int_1__2_), .B(sll_78_ML_int_1__0_), 
        .S(N518), .Z(sll_78_ML_int_2__2_) );
  MUX2_X1 sll_78_M1_1_3 ( .A(sll_78_ML_int_1__3_), .B(sll_78_ML_int_1__1_), 
        .S(N518), .Z(sll_78_ML_int_2__3_) );
  MUX2_X1 sll_78_M1_1_4 ( .A(sll_78_ML_int_1__4_), .B(sll_78_ML_int_1__2_), 
        .S(N518), .Z(sll_78_ML_int_2__4_) );
  MUX2_X1 sll_78_M1_1_5 ( .A(sll_78_ML_int_1__5_), .B(sll_78_ML_int_1__3_), 
        .S(N518), .Z(sll_78_ML_int_2__5_) );
  MUX2_X1 sll_78_M1_1_6 ( .A(sll_78_ML_int_1__6_), .B(sll_78_ML_int_1__4_), 
        .S(N518), .Z(sll_78_ML_int_2__6_) );
  MUX2_X1 sll_78_M1_1_7 ( .A(sll_78_ML_int_1__7_), .B(sll_78_ML_int_1__5_), 
        .S(N518), .Z(sll_78_ML_int_2__7_) );
  MUX2_X1 sll_78_M1_1_8 ( .A(sll_78_ML_int_1__8_), .B(sll_78_ML_int_1__6_), 
        .S(N518), .Z(sll_78_ML_int_2__8_) );
  MUX2_X1 sll_78_M1_1_9 ( .A(sll_78_ML_int_1__9_), .B(sll_78_ML_int_1__7_), 
        .S(N518), .Z(sll_78_ML_int_2__9_) );
  MUX2_X1 sll_78_M1_1_10 ( .A(sll_78_ML_int_1__10_), .B(sll_78_ML_int_1__8_), 
        .S(N518), .Z(sll_78_ML_int_2__10_) );
  MUX2_X1 sll_78_M1_1_11 ( .A(sll_78_ML_int_1__11_), .B(sll_78_ML_int_1__9_), 
        .S(N518), .Z(sll_78_ML_int_2__11_) );
  MUX2_X1 sll_78_M1_1_12 ( .A(sll_78_ML_int_1__12_), .B(sll_78_ML_int_1__10_), 
        .S(N518), .Z(sll_78_ML_int_2__12_) );
  MUX2_X1 sll_78_M1_1_13 ( .A(sll_78_ML_int_1__13_), .B(sll_78_ML_int_1__11_), 
        .S(N518), .Z(sll_78_ML_int_2__13_) );
  MUX2_X1 sll_78_M1_1_14 ( .A(sll_78_ML_int_1__14_), .B(sll_78_ML_int_1__12_), 
        .S(N518), .Z(sll_78_ML_int_2__14_) );
  MUX2_X1 sll_78_M1_1_15 ( .A(sll_78_ML_int_1__15_), .B(sll_78_ML_int_1__13_), 
        .S(N518), .Z(sll_78_ML_int_2__15_) );
  MUX2_X1 sll_78_M1_1_16 ( .A(sll_78_ML_int_1__16_), .B(sll_78_ML_int_1__14_), 
        .S(N518), .Z(sll_78_ML_int_2__16_) );
  MUX2_X1 sll_78_M1_1_17 ( .A(sll_78_ML_int_1__17_), .B(sll_78_ML_int_1__15_), 
        .S(N518), .Z(sll_78_ML_int_2__17_) );
  MUX2_X1 sll_78_M1_1_18 ( .A(sll_78_ML_int_1__18_), .B(sll_78_ML_int_1__16_), 
        .S(N518), .Z(sll_78_ML_int_2__18_) );
  MUX2_X1 sll_78_M1_1_19 ( .A(sll_78_ML_int_1__19_), .B(sll_78_ML_int_1__17_), 
        .S(N518), .Z(sll_78_ML_int_2__19_) );
  MUX2_X1 sll_78_M1_1_20 ( .A(sll_78_ML_int_1__20_), .B(sll_78_ML_int_1__18_), 
        .S(N518), .Z(sll_78_ML_int_2__20_) );
  MUX2_X1 sll_78_M1_1_21 ( .A(sll_78_ML_int_1__21_), .B(sll_78_ML_int_1__19_), 
        .S(N518), .Z(sll_78_ML_int_2__21_) );
  MUX2_X1 sll_78_M1_1_22 ( .A(sll_78_ML_int_1__22_), .B(sll_78_ML_int_1__20_), 
        .S(N518), .Z(sll_78_ML_int_2__22_) );
  MUX2_X1 sll_78_M1_2_4 ( .A(sll_78_ML_int_2__4_), .B(sll_78_ML_int_2__0_), 
        .S(n345), .Z(sll_78_ML_int_3__4_) );
  MUX2_X1 sll_78_M1_2_5 ( .A(sll_78_ML_int_2__5_), .B(sll_78_ML_int_2__1_), 
        .S(n345), .Z(sll_78_ML_int_3__5_) );
  MUX2_X1 sll_78_M1_2_6 ( .A(sll_78_ML_int_2__6_), .B(sll_78_ML_int_2__2_), 
        .S(n345), .Z(sll_78_ML_int_3__6_) );
  MUX2_X1 sll_78_M1_2_7 ( .A(sll_78_ML_int_2__7_), .B(sll_78_ML_int_2__3_), 
        .S(N574), .Z(sll_78_ML_int_3__7_) );
  MUX2_X1 sll_78_M1_2_8 ( .A(sll_78_ML_int_2__8_), .B(sll_78_ML_int_2__4_), 
        .S(N574), .Z(sll_78_ML_int_3__8_) );
  MUX2_X1 sll_78_M1_2_9 ( .A(sll_78_ML_int_2__9_), .B(sll_78_ML_int_2__5_), 
        .S(n345), .Z(sll_78_ML_int_3__9_) );
  MUX2_X1 sll_78_M1_2_10 ( .A(sll_78_ML_int_2__10_), .B(sll_78_ML_int_2__6_), 
        .S(n345), .Z(sll_78_ML_int_3__10_) );
  MUX2_X1 sll_78_M1_2_11 ( .A(sll_78_ML_int_2__11_), .B(sll_78_ML_int_2__7_), 
        .S(n345), .Z(sll_78_ML_int_3__11_) );
  MUX2_X1 sll_78_M1_2_12 ( .A(sll_78_ML_int_2__12_), .B(sll_78_ML_int_2__8_), 
        .S(n345), .Z(sll_78_ML_int_3__12_) );
  MUX2_X1 sll_78_M1_2_13 ( .A(sll_78_ML_int_2__13_), .B(sll_78_ML_int_2__9_), 
        .S(n345), .Z(sll_78_ML_int_3__13_) );
  MUX2_X1 sll_78_M1_2_14 ( .A(sll_78_ML_int_2__14_), .B(sll_78_ML_int_2__10_), 
        .S(n345), .Z(sll_78_ML_int_3__14_) );
  MUX2_X1 sll_78_M1_2_15 ( .A(sll_78_ML_int_2__15_), .B(sll_78_ML_int_2__11_), 
        .S(N574), .Z(sll_78_ML_int_3__15_) );
  MUX2_X1 sll_78_M1_2_16 ( .A(sll_78_ML_int_2__16_), .B(sll_78_ML_int_2__12_), 
        .S(n345), .Z(sll_78_ML_int_3__16_) );
  MUX2_X1 sll_78_M1_2_17 ( .A(sll_78_ML_int_2__17_), .B(sll_78_ML_int_2__13_), 
        .S(N574), .Z(sll_78_ML_int_3__17_) );
  MUX2_X1 sll_78_M1_2_18 ( .A(sll_78_ML_int_2__18_), .B(sll_78_ML_int_2__14_), 
        .S(N574), .Z(sll_78_ML_int_3__18_) );
  MUX2_X1 sll_78_M1_2_19 ( .A(sll_78_ML_int_2__19_), .B(sll_78_ML_int_2__15_), 
        .S(N574), .Z(sll_78_ML_int_3__19_) );
  MUX2_X1 sll_78_M1_2_20 ( .A(sll_78_ML_int_2__20_), .B(sll_78_ML_int_2__16_), 
        .S(N574), .Z(sll_78_ML_int_3__20_) );
  MUX2_X1 sll_78_M1_2_21 ( .A(sll_78_ML_int_2__21_), .B(sll_78_ML_int_2__17_), 
        .S(N574), .Z(sll_78_ML_int_3__21_) );
  MUX2_X1 sll_78_M1_2_22 ( .A(sll_78_ML_int_2__22_), .B(sll_78_ML_int_2__18_), 
        .S(N574), .Z(sll_78_ML_int_3__22_) );
  MUX2_X1 sll_78_M1_3_8 ( .A(sll_78_ML_int_3__8_), .B(sll_78_ML_int_3__0_), 
        .S(N575), .Z(sll_78_ML_int_4__8_) );
  MUX2_X1 sll_78_M1_3_9 ( .A(sll_78_ML_int_3__9_), .B(sll_78_ML_int_3__1_), 
        .S(N575), .Z(sll_78_ML_int_4__9_) );
  MUX2_X1 sll_78_M1_3_10 ( .A(sll_78_ML_int_3__10_), .B(sll_78_ML_int_3__2_), 
        .S(N575), .Z(sll_78_ML_int_4__10_) );
  MUX2_X1 sll_78_M1_3_11 ( .A(sll_78_ML_int_3__11_), .B(sll_78_ML_int_3__3_), 
        .S(N575), .Z(sll_78_ML_int_4__11_) );
  MUX2_X1 sll_78_M1_3_12 ( .A(sll_78_ML_int_3__12_), .B(sll_78_ML_int_3__4_), 
        .S(N575), .Z(sll_78_ML_int_4__12_) );
  MUX2_X1 sll_78_M1_3_13 ( .A(sll_78_ML_int_3__13_), .B(sll_78_ML_int_3__5_), 
        .S(N575), .Z(sll_78_ML_int_4__13_) );
  MUX2_X1 sll_78_M1_3_14 ( .A(sll_78_ML_int_3__14_), .B(sll_78_ML_int_3__6_), 
        .S(N575), .Z(sll_78_ML_int_4__14_) );
  MUX2_X1 sll_78_M1_3_15 ( .A(sll_78_ML_int_3__15_), .B(sll_78_ML_int_3__7_), 
        .S(N575), .Z(sll_78_ML_int_4__15_) );
  MUX2_X1 sll_78_M1_3_16 ( .A(sll_78_ML_int_3__16_), .B(sll_78_ML_int_3__8_), 
        .S(N575), .Z(sll_78_ML_int_4__16_) );
  MUX2_X1 sll_78_M1_3_17 ( .A(sll_78_ML_int_3__17_), .B(sll_78_ML_int_3__9_), 
        .S(N575), .Z(sll_78_ML_int_4__17_) );
  MUX2_X1 sll_78_M1_3_18 ( .A(sll_78_ML_int_3__18_), .B(sll_78_ML_int_3__10_), 
        .S(N575), .Z(sll_78_ML_int_4__18_) );
  MUX2_X1 sll_78_M1_3_19 ( .A(sll_78_ML_int_3__19_), .B(sll_78_ML_int_3__11_), 
        .S(N575), .Z(sll_78_ML_int_4__19_) );
  MUX2_X1 sll_78_M1_3_20 ( .A(sll_78_ML_int_3__20_), .B(sll_78_ML_int_3__12_), 
        .S(N575), .Z(sll_78_ML_int_4__20_) );
  MUX2_X1 sll_78_M1_3_21 ( .A(sll_78_ML_int_3__21_), .B(sll_78_ML_int_3__13_), 
        .S(N575), .Z(sll_78_ML_int_4__21_) );
  MUX2_X1 sll_78_M1_3_22 ( .A(sll_78_ML_int_3__22_), .B(sll_78_ML_int_3__14_), 
        .S(N575), .Z(sll_78_ML_int_4__22_) );
  MUX2_X1 sll_78_M1_4_16 ( .A(sll_78_ML_int_4__16_), .B(n5820), .S(N521), .Z(
        sll_78_ML_int_5__16_) );
  MUX2_X1 sll_78_M1_4_17 ( .A(sll_78_ML_int_4__17_), .B(n578), .S(N521), .Z(
        sll_78_ML_int_5__17_) );
  MUX2_X1 sll_78_M1_4_18 ( .A(sll_78_ML_int_4__18_), .B(n5800), .S(N521), .Z(
        sll_78_ML_int_5__18_) );
  MUX2_X1 sll_78_M1_4_19 ( .A(sll_78_ML_int_4__19_), .B(n5760), .S(N521), .Z(
        sll_78_ML_int_5__19_) );
  MUX2_X1 sll_78_M1_4_20 ( .A(sll_78_ML_int_4__20_), .B(n5810), .S(N521), .Z(
        sll_78_ML_int_5__20_) );
  MUX2_X1 sll_78_M1_4_21 ( .A(sll_78_ML_int_4__21_), .B(n577), .S(N521), .Z(
        sll_78_ML_int_5__21_) );
  MUX2_X1 sll_78_M1_4_22 ( .A(sll_78_ML_int_4__22_), .B(n579), .S(N521), .Z(
        sll_78_ML_int_5__22_) );
  DFF_X1 B_reg_reg_21_ ( .D(n495), .CK(clk), .Q(B_reg[21]), .QN(n1430) );
  DFF_X1 B_reg_reg_22_ ( .D(n496), .CK(clk), .Q(B_reg[22]), .QN(n1420) );
  DFF_X1 A_reg_reg_8_ ( .D(n450), .CK(clk), .Q(A_reg[8]), .QN(n1880) );
  DFF_X1 A_reg_reg_6_ ( .D(n448), .CK(clk), .Q(A_reg[6]), .QN(n1900) );
  DFF_X1 A_reg_reg_5_ ( .D(n447), .CK(clk), .Q(A_reg[5]), .QN(n1910) );
  DFF_X1 A_reg_reg_3_ ( .D(n445), .CK(clk), .Q(A_reg[3]), .QN(n1930) );
  DFF_X1 A_reg_reg_2_ ( .D(n444), .CK(clk), .Q(A_reg[2]), .QN(n1940) );
  DFF_X1 B_reg_reg_31_ ( .D(n505), .CK(clk), .Q(B_reg[31]), .QN(n74) );
  DFF_X1 B_reg_reg_30_ ( .D(n504), .CK(clk), .Q(B_reg[30]), .QN(n604) );
  DFF_X1 B_reg_reg_29_ ( .D(n503), .CK(clk), .Q(B_reg[29]), .QN(n1350) );
  DFF_X1 B_reg_reg_28_ ( .D(n502), .CK(clk), .Q(B_reg[28]), .QN(n603) );
  DFF_X1 B_reg_reg_27_ ( .D(n501), .CK(clk), .Q(B_reg[27]), .QN(n602) );
  DFF_X1 B_reg_reg_26_ ( .D(n500), .CK(clk), .Q(B_reg[26]), .QN(n601) );
  DFF_X1 B_reg_reg_25_ ( .D(n499), .CK(clk), .Q(B_reg[25]), .QN(n600) );
  DFF_X1 B_reg_reg_24_ ( .D(n498), .CK(clk), .Q(B_reg[24]), .QN(n599) );
  DFF_X1 B_reg_reg_23_ ( .D(n497), .CK(clk), .Q(B_reg[23]), .QN(n1410) );
  DFF_X1 A_reg_reg_29_ ( .D(n471), .CK(clk), .Q(A_reg[29]), .QN(n596) );
  DFF_X1 A_reg_reg_23_ ( .D(n465), .CK(clk), .Q(A_reg[23]), .QN(n1730) );
  DFF_X1 A_reg_reg_30_ ( .D(n472), .CK(clk), .Q(A_reg[30]), .QN(n597) );
  DFF_X1 A_reg_reg_28_ ( .D(n470), .CK(clk), .Q(A_reg[28]), .QN(n595) );
  DFF_X1 A_reg_reg_27_ ( .D(n469), .CK(clk), .Q(A_reg[27]), .QN(n594) );
  DFF_X1 A_reg_reg_26_ ( .D(n468), .CK(clk), .Q(A_reg[26]), .QN(n593) );
  DFF_X1 A_reg_reg_25_ ( .D(n467), .CK(clk), .Q(A_reg[25]), .QN(n592) );
  DFF_X1 A_reg_reg_24_ ( .D(n466), .CK(clk), .Q(A_reg[24]), .QN(n1720) );
  DFF_X1 B_reg_reg_20_ ( .D(n494), .CK(clk), .Q(B_reg[20]), .QN(n1440) );
  DFF_X1 B_reg_reg_19_ ( .D(n493), .CK(clk), .Q(B_reg[19]), .QN(n1450) );
  DFF_X1 B_reg_reg_18_ ( .D(n492), .CK(clk), .Q(B_reg[18]), .QN(n1460) );
  DFF_X1 B_reg_reg_17_ ( .D(n491), .CK(clk), .Q(B_reg[17]), .QN(n1470) );
  DFF_X1 B_reg_reg_16_ ( .D(n490), .CK(clk), .Q(B_reg[16]), .QN(n1480) );
  DFF_X1 B_reg_reg_15_ ( .D(n489), .CK(clk), .Q(B_reg[15]), .QN(n1490) );
  DFF_X1 B_reg_reg_14_ ( .D(n488), .CK(clk), .Q(B_reg[14]), .QN(n1500) );
  DFF_X1 B_reg_reg_13_ ( .D(n487), .CK(clk), .Q(B_reg[13]), .QN(n1510) );
  DFF_X1 B_reg_reg_12_ ( .D(n486), .CK(clk), .Q(B_reg[12]), .QN(n1520) );
  DFF_X1 B_reg_reg_11_ ( .D(n485), .CK(clk), .Q(B_reg[11]), .QN(n1530) );
  DFF_X1 B_reg_reg_10_ ( .D(n4840), .CK(clk), .Q(B_reg[10]), .QN(n1540) );
  DFF_X1 B_reg_reg_9_ ( .D(n4830), .CK(clk), .Q(B_reg[9]), .QN(n1550) );
  DFF_X1 B_reg_reg_8_ ( .D(n4820), .CK(clk), .Q(B_reg[8]), .QN(n1560) );
  DFF_X1 B_reg_reg_7_ ( .D(n4810), .CK(clk), .Q(B_reg[7]), .QN(n1570) );
  DFF_X1 B_reg_reg_6_ ( .D(n4800), .CK(clk), .Q(B_reg[6]), .QN(n1580) );
  DFF_X1 B_reg_reg_5_ ( .D(n479), .CK(clk), .Q(B_reg[5]), .QN(n1590) );
  DFF_X1 B_reg_reg_4_ ( .D(n478), .CK(clk), .Q(B_reg[4]), .QN(n1600) );
  DFF_X1 B_reg_reg_3_ ( .D(n477), .CK(clk), .Q(B_reg[3]), .QN(n1610) );
  DFF_X1 B_reg_reg_2_ ( .D(n476), .CK(clk), .Q(B_reg[2]), .QN(n1620) );
  DFF_X1 B_reg_reg_1_ ( .D(n475), .CK(clk), .Q(B_reg[1]), .QN(n1630) );
  DFF_X1 B_reg_reg_0_ ( .D(n474), .CK(clk), .Q(B_reg[0]), .QN(n1640) );
  DFF_X1 A_reg_reg_22_ ( .D(n464), .CK(clk), .Q(A_reg[22]), .QN(n1740) );
  DFF_X1 A_reg_reg_21_ ( .D(n463), .CK(clk), .Q(A_reg[21]), .QN(n1750) );
  DFF_X1 A_reg_reg_20_ ( .D(n462), .CK(clk), .Q(A_reg[20]), .QN(n1760) );
  DFF_X1 A_reg_reg_19_ ( .D(n461), .CK(clk), .Q(A_reg[19]), .QN(n1770) );
  DFF_X1 A_reg_reg_18_ ( .D(n460), .CK(clk), .Q(A_reg[18]), .QN(n1780) );
  DFF_X1 A_reg_reg_17_ ( .D(n459), .CK(clk), .Q(A_reg[17]), .QN(n1790) );
  DFF_X1 A_reg_reg_16_ ( .D(n458), .CK(clk), .Q(A_reg[16]), .QN(n1800) );
  DFF_X1 A_reg_reg_15_ ( .D(n457), .CK(clk), .Q(A_reg[15]), .QN(n1810) );
  DFF_X1 A_reg_reg_14_ ( .D(n456), .CK(clk), .Q(A_reg[14]), .QN(n1820) );
  DFF_X1 A_reg_reg_13_ ( .D(n455), .CK(clk), .Q(A_reg[13]), .QN(n1830) );
  DFF_X1 A_reg_reg_12_ ( .D(n454), .CK(clk), .Q(A_reg[12]), .QN(n1840) );
  DFF_X1 A_reg_reg_11_ ( .D(n453), .CK(clk), .Q(A_reg[11]), .QN(n1850) );
  DFF_X1 A_reg_reg_10_ ( .D(n452), .CK(clk), .Q(A_reg[10]), .QN(n1860) );
  DFF_X1 A_reg_reg_9_ ( .D(n451), .CK(clk), .Q(A_reg[9]), .QN(n1870) );
  DFF_X1 A_reg_reg_7_ ( .D(n449), .CK(clk), .Q(A_reg[7]), .QN(n1890) );
  DFF_X1 A_reg_reg_4_ ( .D(n446), .CK(clk), .Q(A_reg[4]), .QN(n1920) );
  DFF_X1 A_reg_reg_1_ ( .D(n443), .CK(clk), .Q(A_reg[1]), .QN(n1950) );
  DFF_X1 A_reg_reg_0_ ( .D(n442), .CK(clk), .Q(A_reg[0]), .QN(n1960) );
  XNOR2_X1 U518 ( .A(n1650), .B(B_reg[31]), .ZN(n254) );
  OAI22_X1 U519 ( .A1(n548), .A2(n746), .B1(n5620), .B2(n1960), .ZN(MA[0]) );
  OAI21_X1 U520 ( .B1(n5500), .B2(n1640), .A(n426), .ZN(MB[0]) );
  NOR2_X1 U521 ( .A1(n723), .A2(n254), .ZN(n258) );
  INV_X1 U522 ( .A(n346), .ZN(N575) );
  AND2_X1 U523 ( .A1(sub_78_B_4_), .A2(N575), .ZN(n506) );
  INV_X1 U524 ( .A(n542), .ZN(n533) );
  INV_X1 U525 ( .A(n5630), .ZN(n548) );
  INV_X1 U526 ( .A(n5620), .ZN(n546) );
  INV_X1 U527 ( .A(n5620), .ZN(n547) );
  INV_X1 U528 ( .A(n5630), .ZN(n5490) );
  INV_X1 U529 ( .A(n5630), .ZN(n5500) );
  INV_X1 U530 ( .A(n5630), .ZN(n5510) );
  NOR3_X1 U531 ( .A1(sll_78_A_17_), .A2(sll_78_A_19_), .A3(sll_78_A_18_), .ZN(
        n367) );
  INV_X1 U532 ( .A(n573), .ZN(n5750) );
  BUF_X1 U533 ( .A(n543), .Z(n542) );
  BUF_X1 U534 ( .A(n540), .Z(n538) );
  BUF_X1 U535 ( .A(n540), .Z(n539) );
  BUF_X1 U536 ( .A(n543), .Z(n541) );
  BUF_X1 U537 ( .A(n543), .Z(n540) );
  BUF_X1 U538 ( .A(n541), .Z(n534) );
  BUF_X1 U539 ( .A(n536), .Z(n537) );
  BUF_X1 U540 ( .A(n540), .Z(n535) );
  BUF_X1 U541 ( .A(n541), .Z(n536) );
  NOR2_X1 U542 ( .A1(sll_78_A_17_), .A2(sll_78_A_16_), .ZN(n384) );
  INV_X1 U543 ( .A(N484), .ZN(n722) );
  AND2_X1 U544 ( .A1(n351), .A2(n722), .ZN(N483) );
  INV_X1 U545 ( .A(N521), .ZN(n5740) );
  AND2_X1 U546 ( .A1(n252), .A2(N236), .ZN(n508) );
  AND2_X1 U547 ( .A1(n252), .A2(N236), .ZN(n507) );
  AND2_X1 U548 ( .A1(n252), .A2(n723), .ZN(n2050) );
  AND2_X1 U549 ( .A1(n252), .A2(n723), .ZN(n513) );
  AND2_X1 U550 ( .A1(n252), .A2(N236), .ZN(n2070) );
  AND2_X1 U551 ( .A1(n252), .A2(n723), .ZN(n514) );
  NAND4_X1 U552 ( .A1(n354), .A2(n355), .A3(n356), .A4(n357), .ZN(N484) );
  NOR2_X1 U553 ( .A1(sll_78_A_16_), .A2(n358), .ZN(n357) );
  NAND4_X1 U554 ( .A1(n368), .A2(n369), .A3(n370), .A4(n371), .ZN(n363) );
  NAND4_X1 U555 ( .A1(n374), .A2(n375), .A3(n376), .A4(n377), .ZN(n353) );
  NAND4_X1 U556 ( .A1(n378), .A2(n379), .A3(n380), .A4(n381), .ZN(n358) );
  NAND4_X1 U557 ( .A1(n359), .A2(n360), .A3(n361), .A4(n362), .ZN(n351) );
  NOR2_X1 U558 ( .A1(sll_78_A_8_), .A2(n363), .ZN(n362) );
  NOR3_X1 U559 ( .A1(n388), .A2(sll_78_A_11_), .A3(sll_78_A_10_), .ZN(n386) );
  AOI211_X1 U560 ( .C1(n389), .C2(n390), .A(sll_78_A_9_), .B(sll_78_A_8_), 
        .ZN(n388) );
  NOR2_X1 U561 ( .A1(sll_78_A_7_), .A2(sll_78_A_6_), .ZN(n389) );
  NAND3_X1 U562 ( .A1(n374), .A2(n375), .A3(n352), .ZN(n390) );
  OAI211_X1 U563 ( .C1(n382), .C2(n383), .A(n381), .B(n378), .ZN(N481) );
  AOI211_X1 U564 ( .C1(n384), .C2(n385), .A(sll_78_A_19_), .B(sll_78_A_18_), 
        .ZN(n382) );
  NAND2_X1 U565 ( .A1(n379), .A2(n380), .ZN(n383) );
  OAI211_X1 U566 ( .C1(n386), .C2(n387), .A(n370), .B(n371), .ZN(n385) );
  BUF_X1 U567 ( .A(n5640), .Z(n5630) );
  OAI21_X1 U568 ( .B1(sll_78_A_22_), .B2(n393), .A(n378), .ZN(N480) );
  AOI21_X1 U569 ( .B1(n394), .B2(n379), .A(sll_78_A_21_), .ZN(n393) );
  OAI21_X1 U570 ( .B1(sll_78_A_18_), .B2(n395), .A(n355), .ZN(n394) );
  AOI21_X1 U571 ( .B1(n396), .B2(n366), .A(sll_78_A_17_), .ZN(n395) );
  BUF_X1 U572 ( .A(n5640), .Z(n5620) );
  INV_X1 U573 ( .A(n359), .ZN(sll_78_A_10_) );
  INV_X1 U574 ( .A(n354), .ZN(sll_78_A_18_) );
  INV_X1 U575 ( .A(n356), .ZN(sll_78_A_17_) );
  INV_X1 U576 ( .A(n361), .ZN(sll_78_A_9_) );
  OAI21_X1 U577 ( .B1(sll_78_A_6_), .B2(n401), .A(n377), .ZN(n400) );
  AOI21_X1 U578 ( .B1(n402), .B2(n374), .A(sll_78_A_5_), .ZN(n401) );
  OAI21_X1 U579 ( .B1(sll_78_A_2_), .B2(n348), .A(n392), .ZN(n402) );
  OAI21_X1 U580 ( .B1(sll_78_A_14_), .B2(n397), .A(n371), .ZN(n396) );
  AOI21_X1 U581 ( .B1(n398), .B2(n368), .A(sll_78_A_13_), .ZN(n397) );
  OAI21_X1 U582 ( .B1(sll_78_A_10_), .B2(n399), .A(n360), .ZN(n398) );
  AOI21_X1 U583 ( .B1(n400), .B2(n373), .A(sll_78_A_9_), .ZN(n399) );
  NAND2_X1 U584 ( .A1(n391), .A2(n392), .ZN(n352) );
  NAND2_X1 U585 ( .A1(n368), .A2(n369), .ZN(n387) );
  INV_X1 U586 ( .A(n360), .ZN(sll_78_A_11_) );
  BUF_X1 U587 ( .A(n5650), .Z(n5560) );
  BUF_X1 U588 ( .A(n5590), .Z(n5550) );
  BUF_X1 U589 ( .A(n5650), .Z(n5580) );
  BUF_X1 U590 ( .A(n5650), .Z(n5570) );
  INV_X1 U591 ( .A(N278), .ZN(n543) );
  INV_X1 U592 ( .A(n373), .ZN(sll_78_A_8_) );
  INV_X1 U593 ( .A(n366), .ZN(sll_78_A_16_) );
  INV_X1 U594 ( .A(n355), .ZN(sll_78_A_19_) );
  INV_X1 U595 ( .A(n376), .ZN(sll_78_A_6_) );
  INV_X1 U596 ( .A(n377), .ZN(sll_78_A_7_) );
  INV_X1 U597 ( .A(n380), .ZN(sll_78_A_21_) );
  INV_X1 U598 ( .A(n370), .ZN(sll_78_A_14_) );
  INV_X1 U599 ( .A(n369), .ZN(sll_78_A_13_) );
  INV_X1 U600 ( .A(n375), .ZN(sll_78_A_5_) );
  NAND2_X1 U601 ( .A1(n353), .A2(n373), .ZN(n372) );
  INV_X1 U602 ( .A(n381), .ZN(sll_78_A_22_) );
  NAND2_X1 U603 ( .A1(n721), .A2(n364), .ZN(N482) );
  OAI211_X1 U604 ( .C1(n365), .C2(n363), .A(n366), .B(n367), .ZN(n364) );
  INV_X1 U605 ( .A(n358), .ZN(n721) );
  NOR4_X1 U606 ( .A1(n372), .A2(sll_78_A_9_), .A3(sll_78_A_11_), .A4(
        sll_78_A_10_), .ZN(n365) );
  INV_X1 U607 ( .A(n391), .ZN(sll_78_A_2_) );
  INV_X1 U608 ( .A(N236), .ZN(n723) );
  BUF_X1 U609 ( .A(n5590), .Z(n5520) );
  BUF_X1 U610 ( .A(n5610), .Z(n5540) );
  BUF_X1 U611 ( .A(n5530), .Z(n5610) );
  BUF_X1 U612 ( .A(n5520), .Z(n5600) );
  BUF_X1 U613 ( .A(n5570), .Z(n5590) );
  INV_X1 U614 ( .A(n371), .ZN(sll_78_A_15_) );
  INV_X1 U615 ( .A(n379), .ZN(sll_78_A_20_) );
  INV_X1 U616 ( .A(n368), .ZN(sll_78_A_12_) );
  INV_X1 U617 ( .A(n374), .ZN(sll_78_A_4_) );
  INV_X1 U618 ( .A(n392), .ZN(sll_78_A_3_) );
  INV_X1 U619 ( .A(n348), .ZN(sll_78_A_1_) );
  BUF_X1 U620 ( .A(n5590), .Z(n5530) );
  INV_X1 U621 ( .A(MB[23]), .ZN(n635) );
  INV_X1 U622 ( .A(n628), .ZN(n675) );
  XNOR2_X1 U623 ( .A(n347), .B(n346), .ZN(N521) );
  AOI22_X1 U624 ( .A1(N319), .A2(n536), .B1(N295), .B2(n533), .ZN(n371) );
  AOI22_X1 U625 ( .A1(N324), .A2(n535), .B1(N300), .B2(n533), .ZN(n379) );
  AOI22_X1 U626 ( .A1(N316), .A2(n537), .B1(N292), .B2(n533), .ZN(n368) );
  AOI22_X1 U627 ( .A1(N308), .A2(n540), .B1(N284), .B2(n533), .ZN(n374) );
  AOI22_X1 U628 ( .A1(N326), .A2(n534), .B1(N302), .B2(n533), .ZN(n381) );
  AOI22_X1 U629 ( .A1(N325), .A2(n534), .B1(N301), .B2(n533), .ZN(n380) );
  AOI22_X1 U630 ( .A1(N311), .A2(n539), .B1(N287), .B2(n533), .ZN(n377) );
  AOI22_X1 U631 ( .A1(N318), .A2(n536), .B1(N294), .B2(n533), .ZN(n370) );
  AOI22_X1 U632 ( .A1(N312), .A2(n539), .B1(N288), .B2(n533), .ZN(n373) );
  AOI22_X1 U633 ( .A1(N320), .A2(n536), .B1(N296), .B2(n533), .ZN(n366) );
  AOI22_X1 U634 ( .A1(N317), .A2(n537), .B1(N293), .B2(n533), .ZN(n369) );
  AOI22_X1 U635 ( .A1(N309), .A2(n540), .B1(N285), .B2(n533), .ZN(n375) );
  AOI22_X1 U636 ( .A1(N307), .A2(n540), .B1(N283), .B2(n533), .ZN(n392) );
  AOI22_X1 U637 ( .A1(N315), .A2(n537), .B1(N291), .B2(N278), .ZN(n360) );
  AOI22_X1 U638 ( .A1(N323), .A2(n535), .B1(N299), .B2(n533), .ZN(n355) );
  AOI22_X1 U639 ( .A1(N305), .A2(n541), .B1(N281), .B2(n533), .ZN(n348) );
  AOI22_X1 U640 ( .A1(N327), .A2(n534), .B1(N303), .B2(n533), .ZN(n378) );
  AOI22_X1 U641 ( .A1(N313), .A2(n538), .B1(N289), .B2(n533), .ZN(n361) );
  AOI22_X1 U642 ( .A1(N310), .A2(n539), .B1(N286), .B2(n533), .ZN(n376) );
  AOI22_X1 U643 ( .A1(N321), .A2(n535), .B1(N297), .B2(n533), .ZN(n356) );
  AOI22_X1 U644 ( .A1(N306), .A2(n541), .B1(N282), .B2(N278), .ZN(n391) );
  AOI22_X1 U645 ( .A1(N314), .A2(n538), .B1(N290), .B2(N278), .ZN(n359) );
  AOI22_X1 U646 ( .A1(N322), .A2(n538), .B1(N298), .B2(n533), .ZN(n354) );
  AND4_X1 U647 ( .A1(n348), .A2(n722), .A3(n349), .A4(n350), .ZN(n342) );
  NOR3_X1 U648 ( .A1(n351), .A2(n352), .A3(n353), .ZN(n350) );
  AND2_X1 U649 ( .A1(n253), .A2(n748), .ZN(n252) );
  NAND2_X1 U650 ( .A1(sub_78_B_4_), .A2(N575), .ZN(sub_78_carry_5_) );
  BUF_X1 U651 ( .A(n2040), .Z(n509) );
  BUF_X1 U652 ( .A(n2040), .Z(n510) );
  BUF_X1 U653 ( .A(n2040), .Z(n511) );
  BUF_X1 U654 ( .A(n2040), .Z(n512) );
  INV_X1 U655 ( .A(n349), .ZN(sll_78_A_0_) );
  BUF_X1 U656 ( .A(n515), .Z(n5170) );
  BUF_X1 U657 ( .A(n515), .Z(n5180) );
  BUF_X1 U658 ( .A(n515), .Z(n519) );
  BUF_X1 U659 ( .A(n516), .Z(n520) );
  BUF_X1 U660 ( .A(n516), .Z(n5210) );
  BUF_X1 U661 ( .A(n523), .Z(n527) );
  BUF_X1 U662 ( .A(n524), .Z(n528) );
  BUF_X1 U663 ( .A(n524), .Z(n529) );
  BUF_X1 U664 ( .A(n523), .Z(n525) );
  BUF_X1 U665 ( .A(n523), .Z(n526) );
  NOR2_X1 U666 ( .A1(n342), .A2(n748), .ZN(N612) );
  AOI222_X1 U667 ( .A1(N586), .A2(n254), .B1(n263), .B2(N207), .C1(N244), .C2(
        n258), .ZN(n262) );
  AOI222_X1 U668 ( .A1(N582), .A2(n254), .B1(n263), .B2(N203), .C1(N240), .C2(
        n258), .ZN(n267) );
  AOI222_X1 U669 ( .A1(N583), .A2(n254), .B1(n263), .B2(N204), .C1(N241), .C2(
        n258), .ZN(n266) );
  AOI222_X1 U670 ( .A1(N584), .A2(n254), .B1(n263), .B2(N205), .C1(N242), .C2(
        n258), .ZN(n265) );
  AOI222_X1 U671 ( .A1(N581), .A2(n254), .B1(n263), .B2(N202), .C1(N239), .C2(
        n258), .ZN(n1980) );
  AOI222_X1 U672 ( .A1(N585), .A2(n254), .B1(n263), .B2(N206), .C1(N243), .C2(
        n258), .ZN(n264) );
  INV_X1 U673 ( .A(sub_78_B_0_), .ZN(N517) );
  INV_X1 U674 ( .A(n626), .ZN(n674) );
  INV_X1 U675 ( .A(MB[22]), .ZN(n636) );
  INV_X1 U676 ( .A(sub_78_B_1_), .ZN(N518) );
  AOI22_X1 U677 ( .A1(N304), .A2(n541), .B1(N280), .B2(N278), .ZN(n349) );
  INV_X1 U678 ( .A(MA[3]), .ZN(n669) );
  INV_X1 U679 ( .A(MA[2]), .ZN(n668) );
  INV_X1 U680 ( .A(MA[5]), .ZN(n672) );
  INV_X1 U681 ( .A(MA[4]), .ZN(n673) );
  INV_X1 U682 ( .A(MA[7]), .ZN(n670) );
  INV_X1 U683 ( .A(MA[6]), .ZN(n671) );
  INV_X1 U684 ( .A(MA[9]), .ZN(n657) );
  INV_X1 U685 ( .A(MA[8]), .ZN(n658) );
  INV_X1 U686 ( .A(MA[15]), .ZN(n661) );
  INV_X1 U687 ( .A(MA[14]), .ZN(n662) );
  INV_X1 U688 ( .A(MA[17]), .ZN(n655) );
  INV_X1 U689 ( .A(MA[16]), .ZN(n656) );
  INV_X1 U690 ( .A(MA[18]), .ZN(n654) );
  INV_X1 U691 ( .A(MA[19]), .ZN(n653) );
  INV_X1 U692 ( .A(MA[21]), .ZN(n659) );
  INV_X1 U693 ( .A(MA[20]), .ZN(n660) );
  INV_X1 U694 ( .A(MA[11]), .ZN(n665) );
  INV_X1 U695 ( .A(MA[10]), .ZN(n666) );
  INV_X1 U696 ( .A(MA[13]), .ZN(n663) );
  INV_X1 U697 ( .A(MA[12]), .ZN(n664) );
  INV_X1 U698 ( .A(MA[1]), .ZN(n667) );
  INV_X1 U699 ( .A(MA[0]), .ZN(n652) );
  AND2_X1 U700 ( .A1(n253), .A2(n254), .ZN(n2040) );
  AOI222_X1 U701 ( .A1(N580), .A2(n254), .B1(n263), .B2(N201), .C1(N238), .C2(
        n258), .ZN(n2010) );
  NOR2_X1 U702 ( .A1(n747), .A2(n255), .ZN(n253) );
  XNOR2_X1 U703 ( .A(n347), .B(n346), .ZN(N576) );
  INV_X1 U704 ( .A(sub_78_B_2_), .ZN(N574) );
  AND2_X1 U705 ( .A1(n259), .A2(n260), .ZN(n255) );
  NOR4_X1 U706 ( .A1(n264), .A2(n265), .A3(n266), .A4(n267), .ZN(n259) );
  NOR4_X1 U707 ( .A1(n1980), .A2(n2010), .A3(n261), .A4(n262), .ZN(n260) );
  INV_X1 U708 ( .A(MB[1]), .ZN(n645) );
  INV_X1 U709 ( .A(MB[10]), .ZN(n644) );
  INV_X1 U710 ( .A(MB[3]), .ZN(n647) );
  INV_X1 U711 ( .A(MB[5]), .ZN(n650) );
  INV_X1 U712 ( .A(MB[7]), .ZN(n648) );
  INV_X1 U713 ( .A(MB[15]), .ZN(n639) );
  INV_X1 U714 ( .A(MB[2]), .ZN(n646) );
  INV_X1 U715 ( .A(MB[4]), .ZN(n651) );
  INV_X1 U716 ( .A(MB[6]), .ZN(n649) );
  INV_X1 U717 ( .A(MB[8]), .ZN(n634) );
  INV_X1 U718 ( .A(MB[14]), .ZN(n640) );
  INV_X1 U719 ( .A(MB[11]), .ZN(n643) );
  INV_X1 U720 ( .A(MB[13]), .ZN(n641) );
  INV_X1 U721 ( .A(MB[12]), .ZN(n642) );
  INV_X1 U722 ( .A(MB[9]), .ZN(n633) );
  INV_X1 U723 ( .A(n572), .ZN(n579) );
  INV_X1 U724 ( .A(n5710), .ZN(n577) );
  INV_X1 U725 ( .A(n5700), .ZN(n5810) );
  INV_X1 U726 ( .A(n5690), .ZN(n5760) );
  INV_X1 U727 ( .A(n5680), .ZN(n5800) );
  INV_X1 U728 ( .A(n5670), .ZN(n578) );
  INV_X1 U729 ( .A(n5660), .ZN(n5820) );
  INV_X1 U730 ( .A(n2030), .ZN(n718) );
  AOI221_X1 U731 ( .B1(n510), .B2(N571), .C1(n513), .C2(N234), .A(n719), .ZN(
        n2030) );
  INV_X1 U732 ( .A(n2060), .ZN(n719) );
  INV_X1 U733 ( .A(n2080), .ZN(n716) );
  AOI221_X1 U734 ( .B1(n509), .B2(N570), .C1(n2050), .C2(N233), .A(n717), .ZN(
        n2080) );
  INV_X1 U735 ( .A(n209), .ZN(n717) );
  INV_X1 U736 ( .A(n210), .ZN(n714) );
  AOI221_X1 U737 ( .B1(n511), .B2(N569), .C1(n514), .C2(N232), .A(n715), .ZN(
        n210) );
  INV_X1 U738 ( .A(n211), .ZN(n715) );
  INV_X1 U739 ( .A(n2120), .ZN(n712) );
  AOI221_X1 U740 ( .B1(n510), .B2(N568), .C1(n513), .C2(N231), .A(n713), .ZN(
        n2120) );
  INV_X1 U741 ( .A(n2130), .ZN(n713) );
  INV_X1 U742 ( .A(n2140), .ZN(n710) );
  AOI221_X1 U743 ( .B1(n512), .B2(N567), .C1(n2050), .C2(N230), .A(n711), .ZN(
        n2140) );
  INV_X1 U744 ( .A(n2150), .ZN(n711) );
  INV_X1 U745 ( .A(n2160), .ZN(n708) );
  AOI221_X1 U746 ( .B1(n511), .B2(N566), .C1(n514), .C2(N229), .A(n709), .ZN(
        n2160) );
  INV_X1 U747 ( .A(n2170), .ZN(n709) );
  INV_X1 U748 ( .A(n2180), .ZN(n706) );
  AOI221_X1 U749 ( .B1(n510), .B2(N565), .C1(n513), .C2(N228), .A(n707), .ZN(
        n2180) );
  INV_X1 U750 ( .A(n2190), .ZN(n707) );
  INV_X1 U751 ( .A(n2200), .ZN(n704) );
  AOI221_X1 U752 ( .B1(n509), .B2(N564), .C1(n2050), .C2(N227), .A(n705), .ZN(
        n2200) );
  INV_X1 U753 ( .A(n2210), .ZN(n705) );
  INV_X1 U754 ( .A(n2220), .ZN(n702) );
  AOI221_X1 U755 ( .B1(n510), .B2(N563), .C1(n514), .C2(N226), .A(n703), .ZN(
        n2220) );
  INV_X1 U756 ( .A(n2230), .ZN(n703) );
  INV_X1 U757 ( .A(n2240), .ZN(n700) );
  AOI221_X1 U758 ( .B1(n509), .B2(N562), .C1(n513), .C2(N225), .A(n701), .ZN(
        n2240) );
  INV_X1 U759 ( .A(n2250), .ZN(n701) );
  INV_X1 U760 ( .A(n2260), .ZN(n698) );
  AOI221_X1 U761 ( .B1(n509), .B2(N561), .C1(n2050), .C2(N224), .A(n699), .ZN(
        n2260) );
  INV_X1 U762 ( .A(n2270), .ZN(n699) );
  INV_X1 U763 ( .A(n2280), .ZN(n696) );
  AOI221_X1 U764 ( .B1(n512), .B2(N560), .C1(n514), .C2(N223), .A(n697), .ZN(
        n2280) );
  INV_X1 U765 ( .A(n2290), .ZN(n697) );
  INV_X1 U766 ( .A(n2300), .ZN(n694) );
  AOI221_X1 U767 ( .B1(n512), .B2(N559), .C1(n513), .C2(N222), .A(n695), .ZN(
        n2300) );
  INV_X1 U768 ( .A(n2310), .ZN(n695) );
  INV_X1 U769 ( .A(n2320), .ZN(n692) );
  AOI221_X1 U770 ( .B1(n511), .B2(N558), .C1(n2050), .C2(N221), .A(n693), .ZN(
        n2320) );
  INV_X1 U771 ( .A(n2330), .ZN(n693) );
  INV_X1 U772 ( .A(n2340), .ZN(n690) );
  AOI221_X1 U773 ( .B1(n512), .B2(N557), .C1(n514), .C2(N220), .A(n691), .ZN(
        n2340) );
  INV_X1 U774 ( .A(n2350), .ZN(n691) );
  INV_X1 U775 ( .A(n2360), .ZN(n688) );
  AOI221_X1 U776 ( .B1(n511), .B2(N556), .C1(n513), .C2(N219), .A(n689), .ZN(
        n2360) );
  INV_X1 U777 ( .A(n237), .ZN(n689) );
  INV_X1 U778 ( .A(n2380), .ZN(n686) );
  AOI221_X1 U779 ( .B1(n510), .B2(N555), .C1(n2050), .C2(N218), .A(n687), .ZN(
        n2380) );
  INV_X1 U780 ( .A(n2390), .ZN(n687) );
  INV_X1 U781 ( .A(n2400), .ZN(n684) );
  AOI221_X1 U782 ( .B1(n509), .B2(N554), .C1(n514), .C2(N217), .A(n685), .ZN(
        n2400) );
  INV_X1 U783 ( .A(n2410), .ZN(n685) );
  INV_X1 U784 ( .A(n2420), .ZN(n682) );
  AOI221_X1 U785 ( .B1(n511), .B2(N553), .C1(n513), .C2(N216), .A(n683), .ZN(
        n2420) );
  INV_X1 U786 ( .A(n2430), .ZN(n683) );
  INV_X1 U787 ( .A(n2440), .ZN(n680) );
  AOI221_X1 U788 ( .B1(n510), .B2(N552), .C1(n2050), .C2(N215), .A(n681), .ZN(
        n2440) );
  INV_X1 U789 ( .A(n2450), .ZN(n681) );
  INV_X1 U790 ( .A(n246), .ZN(n678) );
  AOI221_X1 U791 ( .B1(n512), .B2(N551), .C1(n2050), .C2(N214), .A(n679), .ZN(
        n246) );
  INV_X1 U792 ( .A(n247), .ZN(n679) );
  INV_X1 U793 ( .A(n248), .ZN(n676) );
  AOI221_X1 U794 ( .B1(n511), .B2(N550), .C1(n513), .C2(N213), .A(n677), .ZN(
        n248) );
  INV_X1 U795 ( .A(n249), .ZN(n677) );
  NOR2_X1 U796 ( .A1(n254), .A2(N236), .ZN(n263) );
  OAI21_X1 U797 ( .B1(n5510), .B2(n749), .A(n411), .ZN(MB[23]) );
  INV_X1 U798 ( .A(IBB), .ZN(n749) );
  NAND2_X1 U799 ( .A1(N168), .A2(n547), .ZN(n411) );
  INV_X1 U800 ( .A(n427), .ZN(r145_B_23_) );
  AOI22_X1 U801 ( .A1(n5520), .A2(N200), .B1(IBA), .B2(n546), .ZN(n427) );
  INV_X1 U802 ( .A(MB[17]), .ZN(n631) );
  INV_X1 U803 ( .A(MB[19]), .ZN(n629) );
  INV_X1 U804 ( .A(MB[21]), .ZN(n637) );
  INV_X1 U805 ( .A(MB[16]), .ZN(n632) );
  INV_X1 U806 ( .A(MB[18]), .ZN(n630) );
  INV_X1 U807 ( .A(MB[20]), .ZN(n638) );
  BUF_X1 U808 ( .A(n2000), .Z(n532) );
  BUF_X1 U809 ( .A(n2000), .Z(n530) );
  BUF_X1 U810 ( .A(n2000), .Z(n531) );
  INV_X1 U811 ( .A(n254), .ZN(n748) );
  INV_X1 U812 ( .A(N177), .ZN(n746) );
  AOI21_X1 U813 ( .B1(n342), .B2(MSB[3]), .A(N483), .ZN(n346) );
  NAND2_X1 U814 ( .A1(N145), .A2(n546), .ZN(n426) );
  OAI22_X1 U815 ( .A1(n5490), .A2(n730), .B1(n5580), .B2(n1950), .ZN(MA[1]) );
  INV_X1 U816 ( .A(N178), .ZN(n730) );
  OAI22_X1 U817 ( .A1(n5490), .A2(n728), .B1(n5560), .B2(n1930), .ZN(MA[3]) );
  INV_X1 U818 ( .A(N180), .ZN(n728) );
  OAI22_X1 U819 ( .A1(n5490), .A2(n725), .B1(n5550), .B2(n1910), .ZN(MA[5]) );
  INV_X1 U820 ( .A(N182), .ZN(n725) );
  OAI22_X1 U821 ( .A1(n5500), .A2(n727), .B1(n5560), .B2(n1890), .ZN(MA[7]) );
  INV_X1 U822 ( .A(N184), .ZN(n727) );
  OAI22_X1 U823 ( .A1(n5490), .A2(n731), .B1(n5620), .B2(n1860), .ZN(MA[10])
         );
  INV_X1 U824 ( .A(N187), .ZN(n731) );
  OAI22_X1 U825 ( .A1(n548), .A2(n734), .B1(n5610), .B2(n1830), .ZN(MA[13]) );
  INV_X1 U826 ( .A(N190), .ZN(n734) );
  OAI22_X1 U827 ( .A1(n5490), .A2(n736), .B1(n5600), .B2(n1810), .ZN(MA[15])
         );
  INV_X1 U828 ( .A(N192), .ZN(n736) );
  OAI22_X1 U829 ( .A1(n5500), .A2(n729), .B1(n5560), .B2(n1940), .ZN(MA[2]) );
  INV_X1 U830 ( .A(N179), .ZN(n729) );
  OAI22_X1 U831 ( .A1(n548), .A2(n724), .B1(n5570), .B2(n1920), .ZN(MA[4]) );
  INV_X1 U832 ( .A(N181), .ZN(n724) );
  OAI22_X1 U833 ( .A1(n548), .A2(n726), .B1(n5550), .B2(n1900), .ZN(MA[6]) );
  INV_X1 U834 ( .A(N183), .ZN(n726) );
  OAI22_X1 U835 ( .A1(n5490), .A2(n740), .B1(n5540), .B2(n1880), .ZN(MA[8]) );
  INV_X1 U836 ( .A(N185), .ZN(n740) );
  OAI22_X1 U837 ( .A1(n5490), .A2(n741), .B1(n5540), .B2(n1870), .ZN(MA[9]) );
  INV_X1 U838 ( .A(N186), .ZN(n741) );
  OAI22_X1 U839 ( .A1(n548), .A2(n733), .B1(n5610), .B2(n1840), .ZN(MA[12]) );
  INV_X1 U840 ( .A(N189), .ZN(n733) );
  OAI22_X1 U841 ( .A1(n548), .A2(n735), .B1(n5600), .B2(n1820), .ZN(MA[14]) );
  INV_X1 U842 ( .A(N191), .ZN(n735) );
  AOI222_X1 U843 ( .A1(N587), .A2(n254), .B1(n263), .B2(N208), .C1(N245), .C2(
        n258), .ZN(n261) );
  OAI22_X1 U844 ( .A1(n5500), .A2(n604), .B1(n5580), .B2(n597), .ZN(N208) );
  OAI21_X1 U845 ( .B1(n5510), .B2(n1620), .A(n410), .ZN(MB[2]) );
  NAND2_X1 U846 ( .A1(N147), .A2(n546), .ZN(n410) );
  OAI21_X1 U847 ( .B1(n5510), .B2(n1600), .A(n408), .ZN(MB[4]) );
  NAND2_X1 U848 ( .A1(N149), .A2(n548), .ZN(n408) );
  OAI21_X1 U849 ( .B1(n5500), .B2(n1580), .A(n406), .ZN(MB[6]) );
  NAND2_X1 U850 ( .A1(N151), .A2(n546), .ZN(n406) );
  OAI21_X1 U851 ( .B1(n5500), .B2(n1560), .A(n404), .ZN(MB[8]) );
  NAND2_X1 U852 ( .A1(N153), .A2(n546), .ZN(n404) );
  OAI21_X1 U853 ( .B1(n5510), .B2(n1500), .A(n421), .ZN(MB[14]) );
  NAND2_X1 U854 ( .A1(N159), .A2(n546), .ZN(n421) );
  OAI21_X1 U855 ( .B1(n5510), .B2(n1630), .A(n415), .ZN(MB[1]) );
  NAND2_X1 U856 ( .A1(N146), .A2(n546), .ZN(n415) );
  OAI21_X1 U857 ( .B1(n545), .B2(n1540), .A(n425), .ZN(MB[10]) );
  NAND2_X1 U858 ( .A1(N155), .A2(n546), .ZN(n425) );
  OAI21_X1 U859 ( .B1(n545), .B2(n1520), .A(n423), .ZN(MB[12]) );
  NAND2_X1 U860 ( .A1(N157), .A2(n547), .ZN(n423) );
  OAI21_X1 U861 ( .B1(n5500), .B2(n1610), .A(n409), .ZN(MB[3]) );
  NAND2_X1 U862 ( .A1(N148), .A2(n547), .ZN(n409) );
  OAI21_X1 U863 ( .B1(n5500), .B2(n1590), .A(n407), .ZN(MB[5]) );
  NAND2_X1 U864 ( .A1(N150), .A2(n547), .ZN(n407) );
  OAI21_X1 U865 ( .B1(n5500), .B2(n1570), .A(n405), .ZN(MB[7]) );
  NAND2_X1 U866 ( .A1(N152), .A2(n546), .ZN(n405) );
  OAI21_X1 U867 ( .B1(n5500), .B2(n1550), .A(n403), .ZN(MB[9]) );
  NAND2_X1 U868 ( .A1(N154), .A2(n546), .ZN(n403) );
  OAI21_X1 U869 ( .B1(n5510), .B2(n1490), .A(n420), .ZN(MB[15]) );
  NAND2_X1 U870 ( .A1(N160), .A2(n546), .ZN(n420) );
  OAI21_X1 U871 ( .B1(n545), .B2(n1530), .A(n424), .ZN(MB[11]) );
  NAND2_X1 U872 ( .A1(N156), .A2(n546), .ZN(n424) );
  OAI21_X1 U873 ( .B1(n545), .B2(n1510), .A(n422), .ZN(MB[13]) );
  NAND2_X1 U874 ( .A1(N158), .A2(n547), .ZN(n422) );
  OAI22_X1 U875 ( .A1(n548), .A2(n732), .B1(n5610), .B2(n1850), .ZN(MA[11]) );
  INV_X1 U876 ( .A(N188), .ZN(n732) );
  INV_X1 U877 ( .A(n5830), .ZN(n598) );
  NAND2_X1 U878 ( .A1(n428), .A2(n429), .ZN(IBB) );
  NOR4_X1 U879 ( .A1(B_reg[26]), .A2(B_reg[25]), .A3(B_reg[24]), .A4(B_reg[23]), .ZN(n428) );
  NOR4_X1 U880 ( .A1(B_reg[30]), .A2(B_reg[29]), .A3(B_reg[28]), .A4(B_reg[27]), .ZN(n429) );
  NAND2_X1 U881 ( .A1(n430), .A2(n431), .ZN(IBA) );
  NOR4_X1 U882 ( .A1(A_reg[30]), .A2(A_reg[29]), .A3(A_reg[28]), .A4(A_reg[27]), .ZN(n431) );
  NOR4_X1 U883 ( .A1(A_reg[26]), .A2(A_reg[25]), .A3(A_reg[24]), .A4(A_reg[23]), .ZN(n430) );
  AOI22_X1 U884 ( .A1(N235), .A2(n508), .B1(result[22]), .B2(n530), .ZN(n2060)
         );
  AOI22_X1 U885 ( .A1(N231), .A2(n508), .B1(result[18]), .B2(n530), .ZN(n2150)
         );
  AOI22_X1 U886 ( .A1(N228), .A2(n508), .B1(result[15]), .B2(n530), .ZN(n2210)
         );
  AOI22_X1 U887 ( .A1(N225), .A2(n508), .B1(result[12]), .B2(n530), .ZN(n2270)
         );
  AOI22_X1 U888 ( .A1(N222), .A2(n508), .B1(result[9]), .B2(n531), .ZN(n2330)
         );
  AOI22_X1 U889 ( .A1(N219), .A2(n508), .B1(result[6]), .B2(n531), .ZN(n2390)
         );
  AOI22_X1 U890 ( .A1(N216), .A2(n508), .B1(result[3]), .B2(n531), .ZN(n2450)
         );
  AOI22_X1 U891 ( .A1(N233), .A2(n507), .B1(result[20]), .B2(n530), .ZN(n211)
         );
  AOI22_X1 U892 ( .A1(N230), .A2(n507), .B1(result[17]), .B2(n530), .ZN(n2170)
         );
  AOI22_X1 U893 ( .A1(N227), .A2(n507), .B1(result[14]), .B2(n530), .ZN(n2230)
         );
  AOI22_X1 U894 ( .A1(N224), .A2(n507), .B1(result[11]), .B2(n530), .ZN(n2290)
         );
  AOI22_X1 U895 ( .A1(N221), .A2(n507), .B1(result[8]), .B2(n531), .ZN(n2350)
         );
  AOI22_X1 U896 ( .A1(N218), .A2(n507), .B1(result[5]), .B2(n531), .ZN(n2410)
         );
  AOI22_X1 U897 ( .A1(N215), .A2(n507), .B1(result[2]), .B2(n531), .ZN(n247)
         );
  AOI22_X1 U898 ( .A1(N232), .A2(n2070), .B1(result[19]), .B2(n530), .ZN(n2130) );
  AOI22_X1 U899 ( .A1(N229), .A2(n2070), .B1(result[16]), .B2(n530), .ZN(n2190) );
  AOI22_X1 U900 ( .A1(N226), .A2(n2070), .B1(result[13]), .B2(n530), .ZN(n2250) );
  AOI22_X1 U901 ( .A1(N223), .A2(n2070), .B1(result[10]), .B2(n531), .ZN(n2310) );
  AOI22_X1 U902 ( .A1(N220), .A2(n2070), .B1(result[7]), .B2(n531), .ZN(n237)
         );
  AOI22_X1 U903 ( .A1(N217), .A2(n2070), .B1(result[4]), .B2(n531), .ZN(n2430)
         );
  AOI22_X1 U904 ( .A1(N214), .A2(n2070), .B1(result[1]), .B2(n531), .ZN(n249)
         );
  AOI22_X1 U905 ( .A1(n507), .A2(N234), .B1(result[21]), .B2(n530), .ZN(n209)
         );
  OAI21_X1 U906 ( .B1(n267), .B2(n747), .A(n341), .ZN(n437) );
  NAND2_X1 U907 ( .A1(result[25]), .A2(n532), .ZN(n341) );
  OAI21_X1 U908 ( .B1(n262), .B2(n747), .A(n337), .ZN(n433) );
  NAND2_X1 U909 ( .A1(result[29]), .A2(n532), .ZN(n337) );
  OAI21_X1 U910 ( .B1(n266), .B2(n747), .A(n340), .ZN(n436) );
  NAND2_X1 U911 ( .A1(result[26]), .A2(n532), .ZN(n340) );
  OAI21_X1 U912 ( .B1(n261), .B2(n747), .A(n336), .ZN(n432) );
  NAND2_X1 U913 ( .A1(result[30]), .A2(n532), .ZN(n336) );
  OAI21_X1 U914 ( .B1(n265), .B2(n747), .A(n339), .ZN(n435) );
  NAND2_X1 U915 ( .A1(result[27]), .A2(n532), .ZN(n339) );
  OAI21_X1 U916 ( .B1(n1980), .B2(n747), .A(n1990), .ZN(n438) );
  NAND2_X1 U917 ( .A1(result[24]), .A2(n531), .ZN(n1990) );
  OAI21_X1 U918 ( .B1(n264), .B2(n747), .A(n338), .ZN(n434) );
  NAND2_X1 U919 ( .A1(result[28]), .A2(n532), .ZN(n338) );
  OAI21_X1 U920 ( .B1(n256), .B2(n747), .A(n257), .ZN(n441) );
  NAND2_X1 U921 ( .A1(overFlow), .A2(n532), .ZN(n257) );
  NOR2_X1 U922 ( .A1(n258), .A2(n255), .ZN(n256) );
  INV_X1 U923 ( .A(n343), .ZN(sub_78_B_0_) );
  AOI21_X1 U924 ( .B1(n342), .B2(MSB[0]), .A(N480), .ZN(n343) );
  INV_X1 U925 ( .A(n345), .ZN(sub_78_B_2_) );
  AOI21_X1 U926 ( .B1(n342), .B2(MSB[2]), .A(N482), .ZN(n345) );
  INV_X1 U927 ( .A(n344), .ZN(sub_78_B_1_) );
  AOI21_X1 U928 ( .B1(n342), .B2(MSB[1]), .A(N481), .ZN(n344) );
  INV_X1 U929 ( .A(n347), .ZN(sub_78_B_4_) );
  AOI21_X1 U930 ( .B1(n342), .B2(MSB[4]), .A(N484), .ZN(n347) );
  AND2_X1 U931 ( .A1(A_reg[23]), .A2(n1410), .ZN(n5830) );
  NAND2_X1 U932 ( .A1(n250), .A2(n251), .ZN(n440) );
  AOI22_X1 U933 ( .A1(N213), .A2(n508), .B1(result[0]), .B2(n531), .ZN(n250)
         );
  AOI22_X1 U934 ( .A1(N549), .A2(n509), .B1(N212), .B2(n514), .ZN(n251) );
  OAI22_X1 U935 ( .A1(n548), .A2(n745), .B1(n5590), .B2(n1770), .ZN(MA[19]) );
  INV_X1 U936 ( .A(N196), .ZN(n745) );
  OAI22_X1 U937 ( .A1(n5490), .A2(n738), .B1(n5570), .B2(n1750), .ZN(MA[21])
         );
  INV_X1 U938 ( .A(N198), .ZN(n738) );
  OAI22_X1 U939 ( .A1(n5500), .A2(n742), .B1(n5600), .B2(n1800), .ZN(MA[16])
         );
  INV_X1 U940 ( .A(N193), .ZN(n742) );
  OAI22_X1 U941 ( .A1(n548), .A2(n744), .B1(n5590), .B2(n1780), .ZN(MA[18]) );
  INV_X1 U942 ( .A(N195), .ZN(n744) );
  OAI22_X1 U943 ( .A1(n548), .A2(n737), .B1(n5580), .B2(n1760), .ZN(MA[20]) );
  INV_X1 U944 ( .A(N197), .ZN(n737) );
  OAI21_X1 U945 ( .B1(n5510), .B2(n1480), .A(n419), .ZN(MB[16]) );
  NAND2_X1 U946 ( .A1(N161), .A2(n547), .ZN(n419) );
  OAI21_X1 U947 ( .B1(n5510), .B2(n1460), .A(n417), .ZN(MB[18]) );
  NAND2_X1 U948 ( .A1(N163), .A2(n547), .ZN(n417) );
  OAI21_X1 U949 ( .B1(n5510), .B2(n1440), .A(n414), .ZN(MB[20]) );
  NAND2_X1 U950 ( .A1(N165), .A2(n547), .ZN(n414) );
  OAI21_X1 U951 ( .B1(n5510), .B2(n1470), .A(n418), .ZN(MB[17]) );
  NAND2_X1 U952 ( .A1(N162), .A2(n547), .ZN(n418) );
  OAI21_X1 U953 ( .B1(n5510), .B2(n1450), .A(n416), .ZN(MB[19]) );
  NAND2_X1 U954 ( .A1(N164), .A2(n547), .ZN(n416) );
  OAI21_X1 U955 ( .B1(n5510), .B2(n1430), .A(n413), .ZN(MB[21]) );
  NAND2_X1 U956 ( .A1(N166), .A2(n547), .ZN(n413) );
  OAI22_X1 U957 ( .A1(n548), .A2(n739), .B1(n5570), .B2(n1740), .ZN(MA[22]) );
  INV_X1 U958 ( .A(N199), .ZN(n739) );
  OAI21_X1 U959 ( .B1(n5510), .B2(n1420), .A(n412), .ZN(MB[22]) );
  NAND2_X1 U960 ( .A1(N167), .A2(n547), .ZN(n412) );
  OAI21_X1 U961 ( .B1(n2010), .B2(n747), .A(n2020), .ZN(n439) );
  NAND2_X1 U962 ( .A1(result[23]), .A2(n532), .ZN(n2020) );
  OAI22_X1 U963 ( .A1(n548), .A2(n743), .B1(n5590), .B2(n1790), .ZN(MA[17]) );
  INV_X1 U964 ( .A(N194), .ZN(n743) );
  OAI22_X1 U965 ( .A1(n5500), .A2(n1410), .B1(n5550), .B2(n1730), .ZN(N201) );
  OAI22_X1 U966 ( .A1(n5490), .A2(n599), .B1(n1720), .B2(n5520), .ZN(N202) );
  INV_X1 U967 ( .A(n334), .ZN(n720) );
  AOI22_X1 U968 ( .A1(n532), .A2(result[31]), .B1(n335), .B2(enable), .ZN(n334) );
  OAI22_X1 U969 ( .A1(n74), .A2(n533), .B1(n1650), .B2(n542), .ZN(n335) );
  OAI22_X1 U970 ( .A1(n5490), .A2(n600), .B1(n5530), .B2(n592), .ZN(N203) );
  OAI22_X1 U971 ( .A1(n5490), .A2(n601), .B1(n5540), .B2(n593), .ZN(N204) );
  OAI22_X1 U972 ( .A1(n5500), .A2(n602), .B1(n5530), .B2(n594), .ZN(N205) );
  OAI22_X1 U973 ( .A1(n5490), .A2(n603), .B1(n5520), .B2(n595), .ZN(N206) );
  OAI22_X1 U974 ( .A1(n5490), .A2(n1350), .B1(n5530), .B2(n596), .ZN(N207) );
  INV_X1 U975 ( .A(enable), .ZN(n747) );
  NOR2_X1 U976 ( .A1(reset), .A2(enable), .ZN(n2000) );
  NOR2_X1 U977 ( .A1(n747), .A2(reset), .ZN(n270) );
  OAI21_X1 U978 ( .B1(n1650), .B2(n525), .A(n3010), .ZN(n473) );
  NAND2_X1 U979 ( .A1(A[31]), .A2(n519), .ZN(n3010) );
  OAI21_X1 U980 ( .B1(n528), .B2(n1960), .A(n269), .ZN(n442) );
  NAND2_X1 U981 ( .A1(A[0]), .A2(n5170), .ZN(n269) );
  OAI21_X1 U982 ( .B1(n527), .B2(n1950), .A(n271), .ZN(n443) );
  NAND2_X1 U983 ( .A1(A[1]), .A2(n5170), .ZN(n271) );
  OAI21_X1 U984 ( .B1(n527), .B2(n1920), .A(n274), .ZN(n446) );
  NAND2_X1 U985 ( .A1(A[4]), .A2(n5170), .ZN(n274) );
  OAI21_X1 U986 ( .B1(n527), .B2(n1890), .A(n277), .ZN(n449) );
  NAND2_X1 U987 ( .A1(A[7]), .A2(n5170), .ZN(n277) );
  OAI21_X1 U988 ( .B1(n527), .B2(n1870), .A(n279), .ZN(n451) );
  NAND2_X1 U989 ( .A1(A[9]), .A2(n5170), .ZN(n279) );
  OAI21_X1 U990 ( .B1(n527), .B2(n1860), .A(n2800), .ZN(n452) );
  NAND2_X1 U991 ( .A1(A[10]), .A2(n5170), .ZN(n2800) );
  OAI21_X1 U992 ( .B1(n527), .B2(n1850), .A(n2810), .ZN(n453) );
  NAND2_X1 U993 ( .A1(A[11]), .A2(n5170), .ZN(n2810) );
  OAI21_X1 U994 ( .B1(n527), .B2(n1840), .A(n2820), .ZN(n454) );
  NAND2_X1 U995 ( .A1(A[12]), .A2(n5180), .ZN(n2820) );
  OAI21_X1 U996 ( .B1(n528), .B2(n1830), .A(n2830), .ZN(n455) );
  NAND2_X1 U997 ( .A1(A[13]), .A2(n5180), .ZN(n2830) );
  OAI21_X1 U998 ( .B1(n527), .B2(n1820), .A(n2840), .ZN(n456) );
  NAND2_X1 U999 ( .A1(A[14]), .A2(n5180), .ZN(n2840) );
  OAI21_X1 U1000 ( .B1(n528), .B2(n1810), .A(n2850), .ZN(n457) );
  NAND2_X1 U1001 ( .A1(A[15]), .A2(n5180), .ZN(n2850) );
  OAI21_X1 U1002 ( .B1(n527), .B2(n1800), .A(n2860), .ZN(n458) );
  NAND2_X1 U1003 ( .A1(A[16]), .A2(n5180), .ZN(n2860) );
  OAI21_X1 U1004 ( .B1(n527), .B2(n1790), .A(n2870), .ZN(n459) );
  NAND2_X1 U1005 ( .A1(A[17]), .A2(n5180), .ZN(n2870) );
  OAI21_X1 U1006 ( .B1(n527), .B2(n1780), .A(n2880), .ZN(n460) );
  NAND2_X1 U1007 ( .A1(A[18]), .A2(n5180), .ZN(n2880) );
  OAI21_X1 U1008 ( .B1(n528), .B2(n1770), .A(n2890), .ZN(n461) );
  NAND2_X1 U1009 ( .A1(A[19]), .A2(n5180), .ZN(n2890) );
  OAI21_X1 U1010 ( .B1(n527), .B2(n1760), .A(n2900), .ZN(n462) );
  NAND2_X1 U1011 ( .A1(A[20]), .A2(n5180), .ZN(n2900) );
  OAI21_X1 U1012 ( .B1(n527), .B2(n1750), .A(n2910), .ZN(n463) );
  NAND2_X1 U1013 ( .A1(A[21]), .A2(n5180), .ZN(n2910) );
  OAI21_X1 U1014 ( .B1(n528), .B2(n1740), .A(n2920), .ZN(n464) );
  NAND2_X1 U1015 ( .A1(A[22]), .A2(n5180), .ZN(n2920) );
  OAI21_X1 U1016 ( .B1(n528), .B2(n1640), .A(n3020), .ZN(n474) );
  NAND2_X1 U1017 ( .A1(B[0]), .A2(n519), .ZN(n3020) );
  OAI21_X1 U1018 ( .B1(n528), .B2(n1630), .A(n3030), .ZN(n475) );
  NAND2_X1 U1019 ( .A1(B[1]), .A2(n519), .ZN(n3030) );
  OAI21_X1 U1020 ( .B1(n528), .B2(n1620), .A(n3040), .ZN(n476) );
  NAND2_X1 U1021 ( .A1(B[2]), .A2(n519), .ZN(n3040) );
  OAI21_X1 U1022 ( .B1(n528), .B2(n1610), .A(n3050), .ZN(n477) );
  NAND2_X1 U1023 ( .A1(B[3]), .A2(n519), .ZN(n3050) );
  OAI21_X1 U1024 ( .B1(n528), .B2(n1600), .A(n3060), .ZN(n478) );
  NAND2_X1 U1025 ( .A1(B[4]), .A2(n520), .ZN(n3060) );
  OAI21_X1 U1026 ( .B1(n528), .B2(n1590), .A(n3070), .ZN(n479) );
  NAND2_X1 U1027 ( .A1(B[5]), .A2(n520), .ZN(n3070) );
  OAI21_X1 U1028 ( .B1(n528), .B2(n1580), .A(n3080), .ZN(n4800) );
  NAND2_X1 U1029 ( .A1(B[6]), .A2(n520), .ZN(n3080) );
  OAI21_X1 U1030 ( .B1(n528), .B2(n1570), .A(n3090), .ZN(n4810) );
  NAND2_X1 U1031 ( .A1(B[7]), .A2(n520), .ZN(n3090) );
  OAI21_X1 U1032 ( .B1(n529), .B2(n1560), .A(n3100), .ZN(n4820) );
  NAND2_X1 U1033 ( .A1(B[8]), .A2(n520), .ZN(n3100) );
  OAI21_X1 U1034 ( .B1(n529), .B2(n1550), .A(n3110), .ZN(n4830) );
  NAND2_X1 U1035 ( .A1(B[9]), .A2(n520), .ZN(n3110) );
  OAI21_X1 U1036 ( .B1(n529), .B2(n1540), .A(n3120), .ZN(n4840) );
  NAND2_X1 U1037 ( .A1(B[10]), .A2(n520), .ZN(n3120) );
  OAI21_X1 U1038 ( .B1(n529), .B2(n1530), .A(n3130), .ZN(n485) );
  NAND2_X1 U1039 ( .A1(B[11]), .A2(n520), .ZN(n3130) );
  OAI21_X1 U1040 ( .B1(n529), .B2(n1520), .A(n3140), .ZN(n486) );
  NAND2_X1 U1041 ( .A1(B[12]), .A2(n520), .ZN(n3140) );
  OAI21_X1 U1042 ( .B1(n529), .B2(n1510), .A(n3150), .ZN(n487) );
  NAND2_X1 U1043 ( .A1(B[13]), .A2(n520), .ZN(n3150) );
  OAI21_X1 U1044 ( .B1(n529), .B2(n1500), .A(n3160), .ZN(n488) );
  NAND2_X1 U1045 ( .A1(B[14]), .A2(n520), .ZN(n3160) );
  OAI21_X1 U1046 ( .B1(n529), .B2(n1490), .A(n3170), .ZN(n489) );
  NAND2_X1 U1047 ( .A1(B[15]), .A2(n520), .ZN(n3170) );
  OAI21_X1 U1048 ( .B1(n529), .B2(n1480), .A(n3180), .ZN(n490) );
  NAND2_X1 U1049 ( .A1(B[16]), .A2(n5210), .ZN(n3180) );
  OAI21_X1 U1050 ( .B1(n529), .B2(n1470), .A(n3190), .ZN(n491) );
  NAND2_X1 U1051 ( .A1(B[17]), .A2(n5210), .ZN(n3190) );
  OAI21_X1 U1052 ( .B1(n529), .B2(n1460), .A(n3200), .ZN(n492) );
  NAND2_X1 U1053 ( .A1(B[18]), .A2(n5210), .ZN(n3200) );
  OAI21_X1 U1054 ( .B1(n529), .B2(n1450), .A(n3210), .ZN(n493) );
  NAND2_X1 U1055 ( .A1(B[19]), .A2(n5210), .ZN(n3210) );
  OAI21_X1 U1056 ( .B1(n529), .B2(n1440), .A(n3220), .ZN(n494) );
  NAND2_X1 U1057 ( .A1(B[20]), .A2(n5210), .ZN(n3220) );
  OAI21_X1 U1058 ( .B1(n1410), .B2(n525), .A(n3250), .ZN(n497) );
  NAND2_X1 U1059 ( .A1(B[23]), .A2(n5210), .ZN(n3250) );
  OAI21_X1 U1060 ( .B1(n599), .B2(n525), .A(n3260), .ZN(n498) );
  NAND2_X1 U1061 ( .A1(B[24]), .A2(n5210), .ZN(n3260) );
  OAI21_X1 U1062 ( .B1(n600), .B2(n525), .A(n3270), .ZN(n499) );
  NAND2_X1 U1063 ( .A1(B[25]), .A2(n5210), .ZN(n3270) );
  OAI21_X1 U1064 ( .B1(n601), .B2(n525), .A(n328), .ZN(n500) );
  NAND2_X1 U1065 ( .A1(B[26]), .A2(n5210), .ZN(n328) );
  OAI21_X1 U1066 ( .B1(n602), .B2(n525), .A(n329), .ZN(n501) );
  NAND2_X1 U1067 ( .A1(B[27]), .A2(n5210), .ZN(n329) );
  OAI21_X1 U1068 ( .B1(n603), .B2(n525), .A(n330), .ZN(n502) );
  NAND2_X1 U1069 ( .A1(B[28]), .A2(n522), .ZN(n330) );
  OAI21_X1 U1070 ( .B1(n1350), .B2(n525), .A(n331), .ZN(n503) );
  NAND2_X1 U1071 ( .A1(B[29]), .A2(n522), .ZN(n331) );
  OAI21_X1 U1072 ( .B1(n604), .B2(n525), .A(n332), .ZN(n504) );
  NAND2_X1 U1073 ( .A1(B[30]), .A2(n522), .ZN(n332) );
  OAI21_X1 U1074 ( .B1(n1730), .B2(n525), .A(n2930), .ZN(n465) );
  NAND2_X1 U1075 ( .A1(A[23]), .A2(n5180), .ZN(n2930) );
  OAI21_X1 U1076 ( .B1(n592), .B2(n526), .A(n2950), .ZN(n467) );
  NAND2_X1 U1077 ( .A1(A[25]), .A2(n519), .ZN(n2950) );
  OAI21_X1 U1078 ( .B1(n593), .B2(n526), .A(n2960), .ZN(n468) );
  NAND2_X1 U1079 ( .A1(A[26]), .A2(n519), .ZN(n2960) );
  OAI21_X1 U1080 ( .B1(n594), .B2(n526), .A(n2970), .ZN(n469) );
  NAND2_X1 U1081 ( .A1(A[27]), .A2(n519), .ZN(n2970) );
  OAI21_X1 U1082 ( .B1(n595), .B2(n526), .A(n2980), .ZN(n470) );
  NAND2_X1 U1083 ( .A1(A[28]), .A2(n519), .ZN(n2980) );
  OAI21_X1 U1084 ( .B1(n596), .B2(n525), .A(n2990), .ZN(n471) );
  NAND2_X1 U1085 ( .A1(A[29]), .A2(n519), .ZN(n2990) );
  OAI21_X1 U1086 ( .B1(n597), .B2(n526), .A(n3000), .ZN(n472) );
  NAND2_X1 U1087 ( .A1(A[30]), .A2(n519), .ZN(n3000) );
  OAI21_X1 U1088 ( .B1(n1720), .B2(n526), .A(n2940), .ZN(n466) );
  NAND2_X1 U1089 ( .A1(A[24]), .A2(n519), .ZN(n2940) );
  OAI21_X1 U1090 ( .B1(n74), .B2(n525), .A(n333), .ZN(n505) );
  NAND2_X1 U1091 ( .A1(B[31]), .A2(n522), .ZN(n333) );
  OAI21_X1 U1092 ( .B1(n526), .B2(n1940), .A(n272), .ZN(n444) );
  NAND2_X1 U1093 ( .A1(A[2]), .A2(n5170), .ZN(n272) );
  OAI21_X1 U1094 ( .B1(n526), .B2(n1930), .A(n273), .ZN(n445) );
  NAND2_X1 U1095 ( .A1(A[3]), .A2(n5170), .ZN(n273) );
  OAI21_X1 U1096 ( .B1(n526), .B2(n1910), .A(n275), .ZN(n447) );
  NAND2_X1 U1097 ( .A1(A[5]), .A2(n5170), .ZN(n275) );
  OAI21_X1 U1098 ( .B1(n526), .B2(n1900), .A(n276), .ZN(n448) );
  NAND2_X1 U1099 ( .A1(A[6]), .A2(n5170), .ZN(n276) );
  OAI21_X1 U1100 ( .B1(n526), .B2(n1880), .A(n2780), .ZN(n450) );
  NAND2_X1 U1101 ( .A1(A[8]), .A2(n5170), .ZN(n2780) );
  OAI21_X1 U1102 ( .B1(n526), .B2(n1420), .A(n3240), .ZN(n496) );
  NAND2_X1 U1103 ( .A1(B[22]), .A2(n5210), .ZN(n3240) );
  OAI21_X1 U1104 ( .B1(n525), .B2(n1430), .A(n3230), .ZN(n495) );
  NAND2_X1 U1105 ( .A1(B[21]), .A2(n5210), .ZN(n3230) );
  OR2_X1 U1106 ( .A1(reset), .A2(n522), .ZN(n268) );
  BUF_X1 U1107 ( .A(n270), .Z(n515) );
  BUF_X1 U1108 ( .A(n270), .Z(n516) );
  BUF_X1 U1109 ( .A(n516), .Z(n522) );
  BUF_X1 U1110 ( .A(n268), .Z(n523) );
  BUF_X1 U1111 ( .A(n268), .Z(n524) );
  BUF_X1 U1112 ( .A(N135), .Z(n544) );
  BUF_X1 U1113 ( .A(N135), .Z(n545) );
  INV_X1 U1114 ( .A(n544), .ZN(n5640) );
  INV_X1 U1115 ( .A(n545), .ZN(n5650) );
  AND2_X1 U1116 ( .A1(sll_78_A_0_), .A2(sub_78_B_0_), .ZN(sll_78_ML_int_1__0_)
         );
  AND2_X1 U1117 ( .A1(sll_78_ML_int_1__0_), .A2(sub_78_B_1_), .ZN(
        sll_78_ML_int_2__0_) );
  AND2_X1 U1118 ( .A1(sll_78_ML_int_1__1_), .A2(sub_78_B_1_), .ZN(
        sll_78_ML_int_2__1_) );
  AND2_X1 U1119 ( .A1(sll_78_ML_int_2__0_), .A2(sub_78_B_2_), .ZN(
        sll_78_ML_int_3__0_) );
  AND2_X1 U1120 ( .A1(sll_78_ML_int_2__1_), .A2(sub_78_B_2_), .ZN(
        sll_78_ML_int_3__1_) );
  AND2_X1 U1121 ( .A1(sll_78_ML_int_2__2_), .A2(sub_78_B_2_), .ZN(
        sll_78_ML_int_3__2_) );
  AND2_X1 U1122 ( .A1(sll_78_ML_int_2__3_), .A2(sub_78_B_2_), .ZN(
        sll_78_ML_int_3__3_) );
  NAND2_X1 U1123 ( .A1(sll_78_ML_int_3__0_), .A2(n346), .ZN(n5660) );
  NAND2_X1 U1124 ( .A1(sll_78_ML_int_3__1_), .A2(n346), .ZN(n5670) );
  NAND2_X1 U1125 ( .A1(sll_78_ML_int_3__2_), .A2(n346), .ZN(n5680) );
  NAND2_X1 U1126 ( .A1(sll_78_ML_int_3__3_), .A2(n346), .ZN(n5690) );
  NAND2_X1 U1127 ( .A1(sll_78_ML_int_3__4_), .A2(n346), .ZN(n5700) );
  NAND2_X1 U1128 ( .A1(sll_78_ML_int_3__5_), .A2(n346), .ZN(n5710) );
  NAND2_X1 U1129 ( .A1(sll_78_ML_int_3__6_), .A2(n346), .ZN(n572) );
  NAND2_X1 U1130 ( .A1(n5740), .A2(sub_78_carry_5_), .ZN(n573) );
  NOR2_X1 U1131 ( .A1(n573), .A2(n5660), .ZN(N549) );
  AND2_X1 U1132 ( .A1(sll_78_ML_int_4__10_), .A2(n5750), .ZN(N559) );
  AND2_X1 U1133 ( .A1(sll_78_ML_int_4__11_), .A2(n5750), .ZN(N560) );
  AND2_X1 U1134 ( .A1(sll_78_ML_int_4__12_), .A2(n5750), .ZN(N561) );
  AND2_X1 U1135 ( .A1(sll_78_ML_int_4__13_), .A2(n5750), .ZN(N562) );
  AND2_X1 U1136 ( .A1(sll_78_ML_int_4__14_), .A2(n5750), .ZN(N563) );
  AND2_X1 U1137 ( .A1(sll_78_ML_int_4__15_), .A2(n5750), .ZN(N564) );
  AND2_X1 U1138 ( .A1(sll_78_ML_int_5__16_), .A2(sub_78_carry_5_), .ZN(N565)
         );
  AND2_X1 U1139 ( .A1(sll_78_ML_int_5__17_), .A2(sub_78_carry_5_), .ZN(N566)
         );
  AND2_X1 U1140 ( .A1(sll_78_ML_int_5__18_), .A2(sub_78_carry_5_), .ZN(N567)
         );
  AND2_X1 U1141 ( .A1(sll_78_ML_int_5__19_), .A2(sub_78_carry_5_), .ZN(N568)
         );
  NOR2_X1 U1142 ( .A1(n573), .A2(n5670), .ZN(N550) );
  AND2_X1 U1143 ( .A1(sll_78_ML_int_5__20_), .A2(sub_78_carry_5_), .ZN(N569)
         );
  AND2_X1 U1144 ( .A1(sll_78_ML_int_5__21_), .A2(sub_78_carry_5_), .ZN(N570)
         );
  AND2_X1 U1145 ( .A1(sll_78_ML_int_5__22_), .A2(sub_78_carry_5_), .ZN(N571)
         );
  NOR2_X1 U1146 ( .A1(n573), .A2(n5680), .ZN(N551) );
  NOR2_X1 U1147 ( .A1(n573), .A2(n5690), .ZN(N552) );
  NOR2_X1 U1148 ( .A1(n573), .A2(n5700), .ZN(N553) );
  NOR2_X1 U1149 ( .A1(n573), .A2(n5710), .ZN(N554) );
  NOR2_X1 U1150 ( .A1(n573), .A2(n572), .ZN(N555) );
  AND3_X1 U1151 ( .A1(n5750), .A2(n346), .A3(sll_78_ML_int_3__7_), .ZN(N556)
         );
  AND2_X1 U1152 ( .A1(sll_78_ML_int_4__8_), .A2(n5750), .ZN(N557) );
  AND2_X1 U1153 ( .A1(sll_78_ML_int_4__9_), .A2(n5750), .ZN(N558) );
  NOR2_X1 U1154 ( .A1(B_reg[29]), .A2(n596), .ZN(n590) );
  AOI21_X1 U1155 ( .B1(n5830), .B2(n599), .A(A_reg[24]), .ZN(n5840) );
  AOI221_X1 U1156 ( .B1(B_reg[25]), .B2(n592), .C1(B_reg[24]), .C2(n598), .A(
        n5840), .ZN(n5850) );
  AOI221_X1 U1157 ( .B1(A_reg[26]), .B2(n601), .C1(A_reg[25]), .C2(n600), .A(
        n5850), .ZN(n5860) );
  AOI221_X1 U1158 ( .B1(B_reg[27]), .B2(n594), .C1(B_reg[26]), .C2(n593), .A(
        n5860), .ZN(n5870) );
  AOI221_X1 U1159 ( .B1(A_reg[28]), .B2(n603), .C1(A_reg[27]), .C2(n602), .A(
        n5870), .ZN(n588) );
  AOI221_X1 U1160 ( .B1(B_reg[29]), .B2(n596), .C1(B_reg[28]), .C2(n595), .A(
        n588), .ZN(n589) );
  OAI22_X1 U1161 ( .A1(n590), .A2(n589), .B1(A_reg[30]), .B2(n604), .ZN(n591)
         );
  OAI21_X1 U1162 ( .B1(B_reg[30]), .B2(n597), .A(n591), .ZN(N135) );
  OAI211_X1 U1163 ( .C1(MB[1]), .C2(n667), .A(n652), .B(MB[0]), .ZN(n605) );
  OAI221_X1 U1164 ( .B1(MA[1]), .B2(n645), .C1(MA[2]), .C2(n646), .A(n605), 
        .ZN(n606) );
  OAI221_X1 U1165 ( .B1(MB[2]), .B2(n668), .C1(MB[3]), .C2(n669), .A(n606), 
        .ZN(n607) );
  OAI221_X1 U1166 ( .B1(MA[3]), .B2(n647), .C1(MA[4]), .C2(n651), .A(n607), 
        .ZN(n608) );
  OAI221_X1 U1167 ( .B1(MB[4]), .B2(n673), .C1(MB[5]), .C2(n672), .A(n608), 
        .ZN(n609) );
  OAI221_X1 U1168 ( .B1(MA[5]), .B2(n650), .C1(MA[6]), .C2(n649), .A(n609), 
        .ZN(n610) );
  OAI221_X1 U1169 ( .B1(MB[6]), .B2(n671), .C1(MB[7]), .C2(n670), .A(n610), 
        .ZN(n611) );
  OAI221_X1 U1170 ( .B1(MA[7]), .B2(n648), .C1(MA[8]), .C2(n634), .A(n611), 
        .ZN(n6120) );
  OAI221_X1 U1171 ( .B1(MB[8]), .B2(n658), .C1(MB[9]), .C2(n657), .A(n6120), 
        .ZN(n613) );
  OAI221_X1 U1172 ( .B1(MA[10]), .B2(n644), .C1(MA[9]), .C2(n633), .A(n613), 
        .ZN(n614) );
  OAI221_X1 U1173 ( .B1(MB[10]), .B2(n666), .C1(MB[11]), .C2(n665), .A(n614), 
        .ZN(n615) );
  OAI221_X1 U1174 ( .B1(MA[11]), .B2(n643), .C1(MA[12]), .C2(n642), .A(n615), 
        .ZN(n616) );
  OAI221_X1 U1175 ( .B1(MB[12]), .B2(n664), .C1(MB[13]), .C2(n663), .A(n616), 
        .ZN(n617) );
  OAI221_X1 U1176 ( .B1(MA[13]), .B2(n641), .C1(MA[14]), .C2(n640), .A(n617), 
        .ZN(n618) );
  OAI221_X1 U1177 ( .B1(MB[14]), .B2(n662), .C1(MB[15]), .C2(n661), .A(n618), 
        .ZN(n619) );
  OAI221_X1 U1178 ( .B1(MA[15]), .B2(n639), .C1(MA[16]), .C2(n632), .A(n619), 
        .ZN(n620) );
  OAI221_X1 U1179 ( .B1(MB[16]), .B2(n656), .C1(MB[17]), .C2(n655), .A(n620), 
        .ZN(n621) );
  OAI221_X1 U1180 ( .B1(MA[17]), .B2(n631), .C1(MA[18]), .C2(n630), .A(n621), 
        .ZN(n622) );
  OAI221_X1 U1181 ( .B1(MB[18]), .B2(n654), .C1(MB[19]), .C2(n653), .A(n622), 
        .ZN(n623) );
  OAI221_X1 U1182 ( .B1(MA[19]), .B2(n629), .C1(MA[20]), .C2(n638), .A(n623), 
        .ZN(n624) );
  OAI221_X1 U1183 ( .B1(MB[20]), .B2(n660), .C1(MB[21]), .C2(n659), .A(n624), 
        .ZN(n625) );
  OAI221_X1 U1184 ( .B1(MA[21]), .B2(n637), .C1(MA[22]), .C2(n636), .A(n625), 
        .ZN(n626) );
  AOI21_X1 U1185 ( .B1(n636), .B2(MA[22]), .A(n674), .ZN(n628) );
  OAI21_X1 U1186 ( .B1(n675), .B2(n635), .A(r145_B_23_), .ZN(n627) );
  OAI21_X1 U1187 ( .B1(MB[23]), .B2(n628), .A(n627), .ZN(N278) );
endmodule

