
module fpAdder_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75;
  wire   [23:1] carry;

  FA_X1 U2_22 ( .A(A[22]), .B(n67), .CI(carry[22]), .CO(carry[23]), .S(
        DIFF[22]) );
  FA_X1 U2_19 ( .A(A[19]), .B(n74), .CI(carry[19]), .CO(carry[20]), .S(
        DIFF[19]) );
  FA_X1 U2_16 ( .A(A[16]), .B(n71), .CI(carry[16]), .CO(carry[17]), .S(
        DIFF[16]) );
  FA_X1 U2_14 ( .A(A[14]), .B(n63), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  FA_X1 U2_13 ( .A(A[13]), .B(n62), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  FA_X1 U2_11 ( .A(A[11]), .B(n60), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  FA_X1 U2_9 ( .A(A[9]), .B(n70), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  FA_X1 U2_7 ( .A(A[7]), .B(n55), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7]) );
  FA_X1 U2_5 ( .A(A[5]), .B(n53), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  FA_X1 U2_4 ( .A(A[4]), .B(n52), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  FA_X1 U2_1 ( .A(A[1]), .B(n58), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  INV_X1 U1 ( .A(B[8]), .ZN(n69) );
  INV_X1 U2 ( .A(B[10]), .ZN(n59) );
  XOR2_X1 U3 ( .A(n66), .B(A[21]), .Z(n1) );
  XOR2_X1 U4 ( .A(n10), .B(n1), .Z(DIFF[21]) );
  NAND2_X1 U5 ( .A1(n9), .A2(n66), .ZN(n2) );
  NAND2_X1 U6 ( .A1(carry[21]), .A2(A[21]), .ZN(n3) );
  NAND2_X1 U7 ( .A1(n66), .A2(A[21]), .ZN(n4) );
  NAND3_X1 U8 ( .A1(n2), .A2(n3), .A3(n4), .ZN(carry[22]) );
  XOR2_X1 U9 ( .A(n59), .B(A[10]), .Z(n5) );
  XOR2_X1 U10 ( .A(carry[10]), .B(n5), .Z(DIFF[10]) );
  NAND2_X1 U11 ( .A1(carry[10]), .A2(n59), .ZN(n6) );
  NAND2_X1 U12 ( .A1(carry[10]), .A2(A[10]), .ZN(n7) );
  NAND2_X1 U13 ( .A1(n59), .A2(A[10]), .ZN(n8) );
  NAND3_X1 U14 ( .A1(n6), .A2(n7), .A3(n8), .ZN(carry[11]) );
  NAND3_X1 U15 ( .A1(n50), .A2(n49), .A3(n51), .ZN(n9) );
  NAND3_X1 U16 ( .A1(n50), .A2(n49), .A3(n51), .ZN(n10) );
  NAND3_X1 U17 ( .A1(n29), .A2(n28), .A3(n30), .ZN(n11) );
  NAND3_X1 U18 ( .A1(n16), .A2(n15), .A3(n17), .ZN(n12) );
  NAND3_X1 U19 ( .A1(n16), .A2(n15), .A3(n17), .ZN(n13) );
  XOR2_X1 U20 ( .A(n57), .B(A[2]), .Z(n14) );
  XOR2_X1 U21 ( .A(carry[2]), .B(n14), .Z(DIFF[2]) );
  NAND2_X1 U22 ( .A1(carry[2]), .A2(n57), .ZN(n15) );
  NAND2_X1 U23 ( .A1(carry[2]), .A2(A[2]), .ZN(n16) );
  NAND2_X1 U24 ( .A1(n57), .A2(A[2]), .ZN(n17) );
  XOR2_X1 U25 ( .A(n56), .B(A[3]), .Z(n18) );
  XOR2_X1 U26 ( .A(n12), .B(n18), .Z(DIFF[3]) );
  NAND2_X1 U27 ( .A1(n13), .A2(n56), .ZN(n19) );
  NAND2_X1 U28 ( .A1(n13), .A2(A[3]), .ZN(n20) );
  NAND2_X1 U29 ( .A1(n56), .A2(A[3]), .ZN(n21) );
  NAND3_X1 U30 ( .A1(n20), .A2(n19), .A3(n21), .ZN(carry[4]) );
  XNOR2_X1 U31 ( .A(carry[23]), .B(n22), .ZN(DIFF[23]) );
  XNOR2_X1 U32 ( .A(A[23]), .B(n68), .ZN(n22) );
  XOR2_X1 U33 ( .A(n69), .B(A[8]), .Z(n23) );
  XOR2_X1 U34 ( .A(carry[8]), .B(n23), .Z(DIFF[8]) );
  NAND2_X1 U35 ( .A1(carry[8]), .A2(n69), .ZN(n24) );
  NAND2_X1 U36 ( .A1(carry[8]), .A2(A[8]), .ZN(n25) );
  NAND2_X1 U37 ( .A1(n69), .A2(A[8]), .ZN(n26) );
  NAND3_X1 U38 ( .A1(n24), .A2(n25), .A3(n26), .ZN(carry[9]) );
  XOR2_X1 U39 ( .A(n72), .B(A[17]), .Z(n27) );
  XOR2_X1 U40 ( .A(carry[17]), .B(n27), .Z(DIFF[17]) );
  NAND2_X1 U41 ( .A1(carry[17]), .A2(n72), .ZN(n28) );
  NAND2_X1 U42 ( .A1(carry[17]), .A2(A[17]), .ZN(n29) );
  NAND2_X1 U43 ( .A1(n72), .A2(A[17]), .ZN(n30) );
  NAND3_X1 U44 ( .A1(n29), .A2(n28), .A3(n30), .ZN(carry[18]) );
  OR2_X1 U45 ( .A1(n75), .A2(A[0]), .ZN(carry[1]) );
  XOR2_X1 U46 ( .A(n61), .B(A[12]), .Z(n31) );
  XOR2_X1 U47 ( .A(carry[12]), .B(n31), .Z(DIFF[12]) );
  NAND2_X1 U48 ( .A1(carry[12]), .A2(n61), .ZN(n32) );
  NAND2_X1 U49 ( .A1(carry[12]), .A2(A[12]), .ZN(n33) );
  NAND2_X1 U50 ( .A1(n61), .A2(A[12]), .ZN(n34) );
  NAND3_X1 U51 ( .A1(n33), .A2(n32), .A3(n34), .ZN(carry[13]) );
  XOR2_X1 U52 ( .A(n54), .B(A[6]), .Z(n35) );
  XOR2_X1 U53 ( .A(carry[6]), .B(n35), .Z(DIFF[6]) );
  NAND2_X1 U54 ( .A1(carry[6]), .A2(n54), .ZN(n36) );
  NAND2_X1 U55 ( .A1(carry[6]), .A2(A[6]), .ZN(n37) );
  NAND2_X1 U56 ( .A1(n54), .A2(A[6]), .ZN(n38) );
  NAND3_X1 U57 ( .A1(n36), .A2(n37), .A3(n38), .ZN(carry[7]) );
  CLKBUF_X1 U58 ( .A(n11), .Z(n39) );
  XOR2_X1 U59 ( .A(n73), .B(A[18]), .Z(n40) );
  XOR2_X1 U60 ( .A(n39), .B(n40), .Z(DIFF[18]) );
  NAND2_X1 U61 ( .A1(carry[18]), .A2(n73), .ZN(n41) );
  NAND2_X1 U62 ( .A1(n11), .A2(A[18]), .ZN(n42) );
  NAND2_X1 U63 ( .A1(n73), .A2(A[18]), .ZN(n43) );
  NAND3_X1 U64 ( .A1(n42), .A2(n41), .A3(n43), .ZN(carry[19]) );
  XOR2_X1 U65 ( .A(n64), .B(A[15]), .Z(n44) );
  XOR2_X1 U66 ( .A(carry[15]), .B(n44), .Z(DIFF[15]) );
  NAND2_X1 U67 ( .A1(carry[15]), .A2(n64), .ZN(n45) );
  NAND2_X1 U68 ( .A1(carry[15]), .A2(A[15]), .ZN(n46) );
  NAND2_X1 U69 ( .A1(n64), .A2(A[15]), .ZN(n47) );
  NAND3_X1 U70 ( .A1(n46), .A2(n45), .A3(n47), .ZN(carry[16]) );
  XOR2_X1 U71 ( .A(n65), .B(A[20]), .Z(n48) );
  XOR2_X1 U72 ( .A(carry[20]), .B(n48), .Z(DIFF[20]) );
  NAND2_X1 U73 ( .A1(carry[20]), .A2(n65), .ZN(n49) );
  NAND2_X1 U74 ( .A1(carry[20]), .A2(A[20]), .ZN(n50) );
  NAND2_X1 U75 ( .A1(n65), .A2(A[20]), .ZN(n51) );
  NAND3_X1 U76 ( .A1(n50), .A2(n49), .A3(n51), .ZN(carry[21]) );
  INV_X1 U77 ( .A(B[23]), .ZN(n68) );
  XNOR2_X1 U78 ( .A(n75), .B(A[0]), .ZN(DIFF[0]) );
  INV_X1 U79 ( .A(B[15]), .ZN(n64) );
  INV_X1 U80 ( .A(B[16]), .ZN(n71) );
  INV_X1 U81 ( .A(B[17]), .ZN(n72) );
  INV_X1 U82 ( .A(B[18]), .ZN(n73) );
  INV_X1 U83 ( .A(B[14]), .ZN(n63) );
  INV_X1 U84 ( .A(B[19]), .ZN(n74) );
  INV_X1 U85 ( .A(B[20]), .ZN(n65) );
  INV_X1 U86 ( .A(B[21]), .ZN(n66) );
  INV_X1 U87 ( .A(B[22]), .ZN(n67) );
  INV_X1 U88 ( .A(B[13]), .ZN(n62) );
  INV_X1 U89 ( .A(B[12]), .ZN(n61) );
  INV_X1 U90 ( .A(B[11]), .ZN(n60) );
  INV_X1 U91 ( .A(B[9]), .ZN(n70) );
  INV_X1 U92 ( .A(B[7]), .ZN(n55) );
  INV_X1 U93 ( .A(B[1]), .ZN(n58) );
  INV_X1 U94 ( .A(B[2]), .ZN(n57) );
  INV_X1 U95 ( .A(B[3]), .ZN(n56) );
  INV_X1 U96 ( .A(B[4]), .ZN(n52) );
  INV_X1 U97 ( .A(B[5]), .ZN(n53) );
  INV_X1 U98 ( .A(B[6]), .ZN(n54) );
  INV_X1 U99 ( .A(B[0]), .ZN(n75) );
endmodule


module fpAdder_DW01_sub_2 ( A, B, CI, DIFF, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81;
  wire   [23:1] carry;

  FA_X1 U2_21 ( .A(A[21]), .B(n72), .CI(carry[21]), .CO(carry[22]), .S(
        DIFF[21]) );
  FA_X1 U2_19 ( .A(A[19]), .B(n80), .CI(carry[19]), .CO(carry[20]), .S(
        DIFF[19]) );
  FA_X1 U2_16 ( .A(A[16]), .B(n77), .CI(carry[16]), .CO(carry[17]), .S(
        DIFF[16]) );
  FA_X1 U2_13 ( .A(A[13]), .B(n68), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  FA_X1 U2_9 ( .A(A[9]), .B(n76), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  FA_X1 U2_7 ( .A(A[7]), .B(n61), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7]) );
  FA_X1 U2_6 ( .A(A[6]), .B(n60), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  FA_X1 U2_4 ( .A(A[4]), .B(n58), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  FA_X1 U2_2 ( .A(A[2]), .B(n63), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  FA_X1 U2_1 ( .A(A[1]), .B(n64), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  XNOR2_X1 U1 ( .A(n74), .B(A[23]), .ZN(n1) );
  CLKBUF_X1 U2 ( .A(n81), .Z(n2) );
  XOR2_X1 U3 ( .A(n73), .B(A[22]), .Z(n3) );
  XOR2_X1 U4 ( .A(carry[22]), .B(n3), .Z(DIFF[22]) );
  NAND2_X1 U5 ( .A1(carry[22]), .A2(n73), .ZN(n4) );
  NAND2_X1 U6 ( .A1(carry[22]), .A2(A[22]), .ZN(n5) );
  NAND2_X1 U7 ( .A1(n73), .A2(A[22]), .ZN(n6) );
  NAND3_X1 U8 ( .A1(n5), .A2(n4), .A3(n6), .ZN(carry[23]) );
  XOR2_X1 U9 ( .A(n59), .B(A[5]), .Z(n7) );
  XOR2_X1 U10 ( .A(carry[5]), .B(n7), .Z(DIFF[5]) );
  NAND2_X1 U11 ( .A1(carry[5]), .A2(n59), .ZN(n8) );
  NAND2_X1 U12 ( .A1(carry[5]), .A2(A[5]), .ZN(n9) );
  NAND2_X1 U13 ( .A1(n59), .A2(A[5]), .ZN(n10) );
  NAND3_X1 U14 ( .A1(n8), .A2(n9), .A3(n10), .ZN(carry[6]) );
  XOR2_X1 U15 ( .A(n71), .B(A[20]), .Z(n11) );
  XOR2_X1 U16 ( .A(carry[20]), .B(n11), .Z(DIFF[20]) );
  NAND2_X1 U17 ( .A1(carry[20]), .A2(n71), .ZN(n12) );
  NAND2_X1 U18 ( .A1(carry[20]), .A2(A[20]), .ZN(n13) );
  NAND2_X1 U19 ( .A1(n71), .A2(A[20]), .ZN(n14) );
  NAND3_X1 U20 ( .A1(n13), .A2(n12), .A3(n14), .ZN(carry[21]) );
  CLKBUF_X1 U21 ( .A(carry[8]), .Z(n15) );
  XOR2_X1 U22 ( .A(n75), .B(A[8]), .Z(n16) );
  XOR2_X1 U23 ( .A(n15), .B(n16), .Z(DIFF[8]) );
  NAND2_X1 U24 ( .A1(carry[8]), .A2(n75), .ZN(n17) );
  NAND2_X1 U25 ( .A1(carry[8]), .A2(A[8]), .ZN(n18) );
  NAND2_X1 U26 ( .A1(n75), .A2(A[8]), .ZN(n19) );
  NAND3_X1 U27 ( .A1(n17), .A2(n18), .A3(n19), .ZN(carry[9]) );
  CLKBUF_X1 U28 ( .A(carry[14]), .Z(n20) );
  XOR2_X1 U29 ( .A(n67), .B(A[12]), .Z(n21) );
  XOR2_X1 U30 ( .A(n25), .B(n21), .Z(DIFF[12]) );
  NAND2_X1 U31 ( .A1(n25), .A2(n67), .ZN(n22) );
  NAND2_X1 U32 ( .A1(carry[12]), .A2(A[12]), .ZN(n23) );
  NAND2_X1 U33 ( .A1(n67), .A2(A[12]), .ZN(n24) );
  NAND3_X1 U34 ( .A1(n22), .A2(n23), .A3(n24), .ZN(carry[13]) );
  NAND3_X1 U35 ( .A1(n31), .A2(n32), .A3(n33), .ZN(n25) );
  XOR2_X1 U36 ( .A(n70), .B(A[15]), .Z(n26) );
  XOR2_X1 U37 ( .A(carry[15]), .B(n26), .Z(DIFF[15]) );
  NAND2_X1 U38 ( .A1(carry[15]), .A2(n70), .ZN(n27) );
  NAND2_X1 U39 ( .A1(carry[15]), .A2(A[15]), .ZN(n28) );
  NAND2_X1 U40 ( .A1(n70), .A2(A[15]), .ZN(n29) );
  NAND3_X1 U41 ( .A1(n28), .A2(n27), .A3(n29), .ZN(carry[16]) );
  XOR2_X1 U42 ( .A(n66), .B(A[11]), .Z(n30) );
  XOR2_X1 U43 ( .A(carry[11]), .B(n30), .Z(DIFF[11]) );
  NAND2_X1 U44 ( .A1(carry[11]), .A2(n66), .ZN(n31) );
  NAND2_X1 U45 ( .A1(carry[11]), .A2(A[11]), .ZN(n32) );
  NAND2_X1 U46 ( .A1(n66), .A2(A[11]), .ZN(n33) );
  NAND3_X1 U47 ( .A1(n31), .A2(n32), .A3(n33), .ZN(carry[12]) );
  CLKBUF_X1 U48 ( .A(n47), .Z(n34) );
  XOR2_X1 U49 ( .A(n79), .B(A[18]), .Z(n35) );
  XOR2_X1 U50 ( .A(n44), .B(n35), .Z(DIFF[18]) );
  NAND2_X1 U51 ( .A1(n43), .A2(n79), .ZN(n36) );
  NAND2_X1 U52 ( .A1(carry[18]), .A2(A[18]), .ZN(n37) );
  NAND2_X1 U53 ( .A1(n79), .A2(A[18]), .ZN(n38) );
  NAND3_X1 U54 ( .A1(n36), .A2(n37), .A3(n38), .ZN(carry[19]) );
  XOR2_X1 U55 ( .A(n69), .B(A[14]), .Z(n39) );
  XOR2_X1 U56 ( .A(n20), .B(n39), .Z(DIFF[14]) );
  NAND2_X1 U57 ( .A1(carry[14]), .A2(n69), .ZN(n40) );
  NAND2_X1 U58 ( .A1(carry[14]), .A2(A[14]), .ZN(n41) );
  NAND2_X1 U59 ( .A1(n69), .A2(A[14]), .ZN(n42) );
  NAND3_X1 U60 ( .A1(n41), .A2(n40), .A3(n42), .ZN(carry[15]) );
  NAND3_X1 U61 ( .A1(n46), .A2(n48), .A3(n47), .ZN(n43) );
  NAND3_X1 U62 ( .A1(n46), .A2(n34), .A3(n48), .ZN(n44) );
  XOR2_X1 U63 ( .A(n78), .B(A[17]), .Z(n45) );
  XOR2_X1 U64 ( .A(carry[17]), .B(n45), .Z(DIFF[17]) );
  NAND2_X1 U65 ( .A1(carry[17]), .A2(n78), .ZN(n46) );
  NAND2_X1 U66 ( .A1(carry[17]), .A2(A[17]), .ZN(n47) );
  NAND2_X1 U67 ( .A1(n78), .A2(A[17]), .ZN(n48) );
  NAND3_X1 U68 ( .A1(n46), .A2(n47), .A3(n48), .ZN(carry[18]) );
  XNOR2_X1 U69 ( .A(carry[23]), .B(n1), .ZN(DIFF[23]) );
  XOR2_X1 U70 ( .A(n62), .B(A[3]), .Z(n49) );
  XOR2_X1 U71 ( .A(carry[3]), .B(n49), .Z(DIFF[3]) );
  NAND2_X1 U72 ( .A1(carry[3]), .A2(n62), .ZN(n50) );
  NAND2_X1 U73 ( .A1(carry[3]), .A2(A[3]), .ZN(n51) );
  NAND2_X1 U74 ( .A1(n62), .A2(A[3]), .ZN(n52) );
  NAND3_X1 U75 ( .A1(n51), .A2(n50), .A3(n52), .ZN(carry[4]) );
  XOR2_X1 U76 ( .A(n65), .B(A[10]), .Z(n53) );
  XOR2_X1 U77 ( .A(carry[10]), .B(n53), .Z(DIFF[10]) );
  NAND2_X1 U78 ( .A1(carry[10]), .A2(n65), .ZN(n54) );
  NAND2_X1 U79 ( .A1(carry[10]), .A2(A[10]), .ZN(n55) );
  NAND2_X1 U80 ( .A1(n65), .A2(A[10]), .ZN(n56) );
  NAND3_X1 U81 ( .A1(n54), .A2(n55), .A3(n56), .ZN(carry[11]) );
  XNOR2_X1 U82 ( .A(A[0]), .B(n2), .ZN(DIFF[0]) );
  INV_X1 U83 ( .A(B[23]), .ZN(n74) );
  INV_X1 U84 ( .A(B[15]), .ZN(n70) );
  INV_X1 U85 ( .A(B[16]), .ZN(n77) );
  INV_X1 U86 ( .A(B[17]), .ZN(n78) );
  INV_X1 U87 ( .A(B[18]), .ZN(n79) );
  INV_X1 U88 ( .A(B[14]), .ZN(n69) );
  INV_X1 U89 ( .A(B[19]), .ZN(n80) );
  INV_X1 U90 ( .A(B[20]), .ZN(n71) );
  INV_X1 U91 ( .A(B[21]), .ZN(n72) );
  INV_X1 U92 ( .A(B[22]), .ZN(n73) );
  INV_X1 U93 ( .A(B[13]), .ZN(n68) );
  INV_X1 U94 ( .A(B[12]), .ZN(n67) );
  INV_X1 U95 ( .A(B[11]), .ZN(n66) );
  INV_X1 U96 ( .A(B[10]), .ZN(n65) );
  INV_X1 U97 ( .A(B[9]), .ZN(n76) );
  INV_X1 U98 ( .A(B[8]), .ZN(n75) );
  INV_X1 U99 ( .A(B[7]), .ZN(n61) );
  INV_X1 U100 ( .A(B[6]), .ZN(n60) );
  INV_X1 U101 ( .A(B[1]), .ZN(n64) );
  NAND2_X1 U102 ( .A1(B[0]), .A2(n57), .ZN(carry[1]) );
  INV_X1 U103 ( .A(A[0]), .ZN(n57) );
  INV_X1 U104 ( .A(B[2]), .ZN(n63) );
  INV_X1 U105 ( .A(B[3]), .ZN(n62) );
  INV_X1 U106 ( .A(B[4]), .ZN(n58) );
  INV_X1 U107 ( .A(B[5]), .ZN(n59) );
  INV_X1 U108 ( .A(B[0]), .ZN(n81) );
endmodule


module fpAdder_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HA_X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  HA_X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  HA_X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  HA_X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  HA_X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  HA_X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  INV_X1 U1 ( .A(A[0]), .ZN(SUM[0]) );
  XOR2_X1 U2 ( .A(carry[7]), .B(A[7]), .Z(SUM[7]) );
endmodule


module fpAdder_DW01_add_0 ( A, B, CI, SUM, CO );
  input [24:0] A;
  input [24:0] B;
  output [24:0] SUM;
  input CI;
  output CO;

  wire   [23:1] carry;

  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(SUM[24]), .S(SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  FA_X1 U1_0 ( .A(A[0]), .B(B[0]), .CI(1'b0), .CO(carry[1]), .S(SUM[0]) );
endmodule


module fpAdder_DW_rash_0 ( A, DATA_TC, SH, SH_TC, B );
  input [23:0] A;
  input [7:0] SH;
  output [23:0] B;
  input DATA_TC, SH_TC;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155;

  NAND2_X1 U3 ( .A1(n111), .A2(n99), .ZN(n1) );
  NAND2_X1 U4 ( .A1(n112), .A2(n98), .ZN(n2) );
  NAND2_X1 U5 ( .A1(n114), .A2(n96), .ZN(n3) );
  AND3_X1 U6 ( .A1(n1), .A2(n2), .A3(n3), .ZN(n149) );
  INV_X1 U7 ( .A(SH[2]), .ZN(n24) );
  OR2_X2 U8 ( .A1(n7), .A2(n12), .ZN(n11) );
  OR2_X1 U9 ( .A1(SH[5]), .A2(SH[3]), .ZN(n12) );
  NOR2_X1 U10 ( .A1(SH[6]), .A2(n12), .ZN(n148) );
  NOR2_X2 U11 ( .A1(n7), .A2(n8), .ZN(n111) );
  OR2_X1 U12 ( .A1(n5), .A2(n73), .ZN(n4) );
  CLKBUF_X1 U13 ( .A(n11), .Z(n5) );
  OR2_X1 U14 ( .A1(SH[5]), .A2(n6), .ZN(n8) );
  OR2_X1 U15 ( .A1(SH[3]), .A2(n24), .ZN(n6) );
  BUF_X1 U16 ( .A(SH[6]), .Z(n7) );
  AOI222_X1 U17 ( .A1(n111), .A2(n86), .B1(n112), .B2(n123), .C1(n114), .C2(
        n84), .ZN(n122) );
  NOR2_X1 U18 ( .A1(SH[4]), .A2(n150), .ZN(n9) );
  NOR2_X1 U19 ( .A1(SH[4]), .A2(n150), .ZN(n10) );
  NAND2_X1 U20 ( .A1(n111), .A2(n22), .ZN(n72) );
  INV_X1 U21 ( .A(n133), .ZN(n22) );
  INV_X1 U22 ( .A(n75), .ZN(n21) );
  INV_X1 U23 ( .A(n80), .ZN(n36) );
  INV_X1 U24 ( .A(n90), .ZN(n39) );
  INV_X1 U25 ( .A(n85), .ZN(n31) );
  INV_X1 U26 ( .A(SH[0]), .ZN(n46) );
  INV_X1 U27 ( .A(n76), .ZN(n34) );
  INV_X1 U28 ( .A(n96), .ZN(n29) );
  INV_X1 U29 ( .A(n89), .ZN(n38) );
  INV_X1 U30 ( .A(n84), .ZN(n33) );
  INV_X1 U31 ( .A(n94), .ZN(n25) );
  INV_X1 U32 ( .A(SH[7]), .ZN(n23) );
  INV_X1 U33 ( .A(n113), .ZN(n35) );
  INV_X1 U34 ( .A(n98), .ZN(n28) );
  INV_X1 U35 ( .A(n91), .ZN(n42) );
  INV_X1 U36 ( .A(n123), .ZN(n30) );
  INV_X1 U37 ( .A(n88), .ZN(n40) );
  INV_X1 U38 ( .A(n95), .ZN(n26) );
  INV_X1 U39 ( .A(n83), .ZN(n32) );
  INV_X1 U40 ( .A(n78), .ZN(n37) );
  INV_X1 U41 ( .A(n105), .ZN(n45) );
  INV_X1 U42 ( .A(n92), .ZN(n41) );
  INV_X1 U43 ( .A(n81), .ZN(n44) );
  INV_X1 U44 ( .A(A[23]), .ZN(n47) );
  INV_X1 U45 ( .A(n99), .ZN(n27) );
  INV_X1 U46 ( .A(n86), .ZN(n43) );
  INV_X1 U47 ( .A(A[2]), .ZN(n68) );
  INV_X1 U48 ( .A(A[22]), .ZN(n48) );
  INV_X1 U49 ( .A(A[21]), .ZN(n49) );
  INV_X1 U50 ( .A(A[20]), .ZN(n50) );
  INV_X1 U51 ( .A(A[19]), .ZN(n51) );
  INV_X1 U52 ( .A(A[18]), .ZN(n52) );
  INV_X1 U53 ( .A(A[11]), .ZN(n59) );
  INV_X1 U54 ( .A(A[10]), .ZN(n60) );
  INV_X1 U55 ( .A(A[14]), .ZN(n56) );
  INV_X1 U56 ( .A(A[15]), .ZN(n55) );
  INV_X1 U57 ( .A(A[6]), .ZN(n64) );
  INV_X1 U58 ( .A(A[7]), .ZN(n63) );
  INV_X1 U59 ( .A(A[16]), .ZN(n54) );
  INV_X1 U60 ( .A(A[3]), .ZN(n67) );
  INV_X1 U61 ( .A(A[12]), .ZN(n58) );
  INV_X1 U62 ( .A(A[4]), .ZN(n66) );
  INV_X1 U63 ( .A(A[13]), .ZN(n57) );
  INV_X1 U64 ( .A(A[5]), .ZN(n65) );
  INV_X1 U65 ( .A(A[8]), .ZN(n62) );
  INV_X1 U66 ( .A(A[17]), .ZN(n53) );
  INV_X1 U67 ( .A(A[9]), .ZN(n61) );
  BUF_X2 U68 ( .A(n108), .Z(n19) );
  BUF_X2 U69 ( .A(n108), .Z(n20) );
  NAND2_X2 U70 ( .A1(n102), .A2(n23), .ZN(n69) );
  NOR2_X1 U71 ( .A1(n46), .A2(SH[1]), .ZN(n13) );
  NOR2_X1 U72 ( .A1(n46), .A2(SH[1]), .ZN(n14) );
  NAND2_X1 U73 ( .A1(n46), .A2(SH[1]), .ZN(n15) );
  NAND2_X1 U74 ( .A1(n46), .A2(SH[1]), .ZN(n16) );
  NAND2_X1 U75 ( .A1(SH[0]), .A2(SH[1]), .ZN(n17) );
  NAND2_X1 U76 ( .A1(SH[0]), .A2(SH[1]), .ZN(n18) );
  OAI222_X1 U77 ( .A1(n42), .A2(n69), .B1(n70), .B2(n71), .C1(n38), .C2(n72), 
        .ZN(B[9]) );
  OAI222_X1 U78 ( .A1(n28), .A2(n69), .B1(n73), .B2(n71), .C1(n29), .C2(n72), 
        .ZN(B[8]) );
  OAI221_X1 U79 ( .B1(n44), .B2(n69), .C1(n35), .C2(n72), .A(n74), .ZN(B[7])
         );
  AOI222_X1 U80 ( .A1(n75), .A2(n76), .B1(n77), .B2(n78), .C1(n79), .C2(n36), 
        .ZN(n74) );
  OAI221_X1 U81 ( .B1(n43), .B2(n69), .C1(n30), .C2(n72), .A(n82), .ZN(B[6])
         );
  AOI222_X1 U82 ( .A1(n79), .A2(n31), .B1(n77), .B2(n83), .C1(n75), .C2(n84), 
        .ZN(n82) );
  OAI221_X1 U83 ( .B1(n41), .B2(n69), .C1(n42), .C2(n72), .A(n87), .ZN(B[5])
         );
  AOI222_X1 U84 ( .A1(n79), .A2(n39), .B1(n77), .B2(n88), .C1(n75), .C2(n89), 
        .ZN(n87) );
  OAI221_X1 U85 ( .B1(n27), .B2(n69), .C1(n28), .C2(n72), .A(n93), .ZN(B[4])
         );
  AOI222_X1 U86 ( .A1(n79), .A2(n94), .B1(n77), .B2(n95), .C1(n75), .C2(n96), 
        .ZN(n93) );
  NOR2_X1 U87 ( .A1(n71), .A2(n24), .ZN(n77) );
  NOR4_X1 U88 ( .A1(n5), .A2(SH[2]), .A3(n10), .A4(SH[7]), .ZN(n79) );
  AOI21_X1 U89 ( .B1(n100), .B2(n101), .A(SH[7]), .ZN(B[3]) );
  NAND2_X1 U90 ( .A1(n102), .A2(n103), .ZN(n101) );
  OAI221_X1 U91 ( .B1(n104), .B2(n64), .C1(n15), .C2(n65), .A(n106), .ZN(n103)
         );
  AOI22_X1 U92 ( .A1(A[4]), .A2(n14), .B1(A[3]), .B2(n19), .ZN(n106) );
  MUX2_X1 U93 ( .A(n109), .B(n110), .S(n9), .Z(n100) );
  AOI222_X1 U94 ( .A1(n111), .A2(n81), .B1(n112), .B2(n113), .C1(n114), .C2(
        n76), .ZN(n110) );
  OAI221_X1 U95 ( .B1(n18), .B2(n60), .C1(n105), .C2(n61), .A(n115), .ZN(n81)
         );
  AOI22_X1 U96 ( .A1(A[8]), .A2(n13), .B1(A[7]), .B2(n19), .ZN(n115) );
  OR2_X1 U97 ( .A1(n5), .A2(n116), .ZN(n109) );
  AOI21_X1 U98 ( .B1(n117), .B2(n118), .A(SH[7]), .ZN(B[2]) );
  NAND2_X1 U99 ( .A1(n102), .A2(n119), .ZN(n118) );
  OAI221_X1 U100 ( .B1(n17), .B2(n65), .C1(n16), .C2(n66), .A(n120), .ZN(n119)
         );
  AOI22_X1 U101 ( .A1(A[3]), .A2(n107), .B1(A[2]), .B2(n19), .ZN(n120) );
  MUX2_X1 U102 ( .A(n121), .B(n122), .S(n10), .Z(n117) );
  OAI221_X1 U103 ( .B1(n104), .B2(n61), .C1(n15), .C2(n62), .A(n124), .ZN(n86)
         );
  AOI22_X1 U104 ( .A1(A[7]), .A2(n14), .B1(A[6]), .B2(n19), .ZN(n124) );
  NOR2_X1 U105 ( .A1(n69), .A2(n80), .ZN(B[23]) );
  NOR2_X1 U106 ( .A1(n85), .A2(n69), .ZN(B[22]) );
  NOR2_X1 U107 ( .A1(n90), .A2(n69), .ZN(B[21]) );
  NOR2_X1 U108 ( .A1(n25), .A2(n69), .ZN(B[20]) );
  AOI21_X1 U109 ( .B1(n125), .B2(n126), .A(SH[7]), .ZN(B[1]) );
  NAND2_X1 U110 ( .A1(n102), .A2(n127), .ZN(n126) );
  OAI221_X1 U111 ( .B1(n18), .B2(n66), .C1(n105), .C2(n67), .A(n128), .ZN(n127) );
  AOI22_X1 U112 ( .A1(A[2]), .A2(n13), .B1(A[1]), .B2(n19), .ZN(n128) );
  MUX2_X1 U113 ( .A(n129), .B(n130), .S(n9), .Z(n125) );
  AOI222_X1 U114 ( .A1(n111), .A2(n92), .B1(n112), .B2(n91), .C1(n114), .C2(
        n89), .ZN(n130) );
  OAI221_X1 U115 ( .B1(n17), .B2(n58), .C1(n16), .C2(n59), .A(n131), .ZN(n91)
         );
  AOI22_X1 U116 ( .A1(A[10]), .A2(n107), .B1(A[9]), .B2(n19), .ZN(n131) );
  OAI221_X1 U117 ( .B1(n104), .B2(n62), .C1(n15), .C2(n63), .A(n132), .ZN(n92)
         );
  AOI22_X1 U118 ( .A1(A[6]), .A2(n14), .B1(A[5]), .B2(n19), .ZN(n132) );
  NOR3_X1 U119 ( .A1(n5), .A2(n116), .A3(n133), .ZN(B[19]) );
  NOR2_X1 U120 ( .A1(n133), .A2(n121), .ZN(B[18]) );
  OR2_X1 U121 ( .A1(n11), .A2(n134), .ZN(n121) );
  NOR2_X1 U122 ( .A1(n133), .A2(n129), .ZN(B[17]) );
  OR2_X1 U123 ( .A1(n11), .A2(n70), .ZN(n129) );
  MUX2_X1 U124 ( .A(n90), .B(n40), .S(n24), .Z(n70) );
  NOR2_X1 U125 ( .A1(n133), .A2(n4), .ZN(B[16]) );
  OAI222_X1 U126 ( .A1(n34), .A2(n69), .B1(n80), .B2(n21), .C1(n37), .C2(n72), 
        .ZN(B[15]) );
  OAI222_X1 U127 ( .A1(n33), .A2(n69), .B1(n85), .B2(n21), .C1(n32), .C2(n72), 
        .ZN(B[14]) );
  OAI222_X1 U128 ( .A1(n38), .A2(n69), .B1(n90), .B2(n21), .C1(n40), .C2(n72), 
        .ZN(B[13]) );
  OAI221_X1 U129 ( .B1(n18), .B2(n50), .C1(n105), .C2(n51), .A(n136), .ZN(n88)
         );
  AOI22_X1 U130 ( .A1(A[18]), .A2(n13), .B1(A[17]), .B2(n19), .ZN(n136) );
  AOI222_X1 U131 ( .A1(n13), .A2(A[22]), .B1(n45), .B2(A[23]), .C1(n20), .C2(
        A[21]), .ZN(n90) );
  OAI221_X1 U132 ( .B1(n17), .B2(n54), .C1(n16), .C2(n55), .A(n137), .ZN(n89)
         );
  AOI22_X1 U133 ( .A1(A[14]), .A2(n107), .B1(A[13]), .B2(n19), .ZN(n137) );
  OAI222_X1 U134 ( .A1(n29), .A2(n69), .B1(n25), .B2(n21), .C1(n26), .C2(n72), 
        .ZN(B[12]) );
  NOR2_X1 U135 ( .A1(n71), .A2(SH[2]), .ZN(n75) );
  OAI222_X1 U136 ( .A1(n34), .A2(n72), .B1(n35), .B2(n69), .C1(n116), .C2(n71), 
        .ZN(B[11]) );
  MUX2_X1 U137 ( .A(n80), .B(n37), .S(n24), .Z(n116) );
  OAI221_X1 U138 ( .B1(n48), .B2(n104), .C1(n15), .C2(n49), .A(n138), .ZN(n78)
         );
  AOI22_X1 U139 ( .A1(A[20]), .A2(n14), .B1(A[19]), .B2(n19), .ZN(n138) );
  NAND2_X1 U140 ( .A1(n20), .A2(A[23]), .ZN(n80) );
  OAI221_X1 U141 ( .B1(n104), .B2(n56), .C1(n105), .C2(n57), .A(n139), .ZN(
        n113) );
  AOI22_X1 U142 ( .A1(A[12]), .A2(n13), .B1(A[11]), .B2(n20), .ZN(n139) );
  OAI221_X1 U143 ( .B1(n18), .B2(n52), .C1(n16), .C2(n53), .A(n140), .ZN(n76)
         );
  AOI22_X1 U144 ( .A1(A[16]), .A2(n107), .B1(A[15]), .B2(n20), .ZN(n140) );
  OAI222_X1 U145 ( .A1(n30), .A2(n69), .B1(n134), .B2(n71), .C1(n33), .C2(n72), 
        .ZN(B[10]) );
  OAI221_X1 U146 ( .B1(n17), .B2(n53), .C1(n15), .C2(n54), .A(n141), .ZN(n84)
         );
  AOI22_X1 U147 ( .A1(A[15]), .A2(n14), .B1(A[14]), .B2(n20), .ZN(n141) );
  NAND2_X1 U148 ( .A1(n22), .A2(n11), .ZN(n71) );
  NAND2_X1 U149 ( .A1(n9), .A2(n23), .ZN(n133) );
  MUX2_X1 U150 ( .A(n85), .B(n32), .S(n24), .Z(n134) );
  OAI221_X1 U151 ( .B1(n49), .B2(n18), .C1(n105), .C2(n50), .A(n142), .ZN(n83)
         );
  AOI22_X1 U152 ( .A1(A[19]), .A2(n13), .B1(A[18]), .B2(n20), .ZN(n142) );
  AOI22_X1 U153 ( .A1(A[22]), .A2(n19), .B1(A[23]), .B2(n14), .ZN(n85) );
  OAI221_X1 U154 ( .B1(n104), .B2(n57), .C1(n16), .C2(n58), .A(n143), .ZN(n123) );
  AOI22_X1 U155 ( .A1(A[11]), .A2(n107), .B1(A[10]), .B2(n20), .ZN(n143) );
  AOI21_X1 U156 ( .B1(n144), .B2(n145), .A(SH[7]), .ZN(B[0]) );
  NAND2_X1 U157 ( .A1(n102), .A2(n146), .ZN(n145) );
  OAI221_X1 U158 ( .B1(n18), .B2(n67), .C1(n15), .C2(n68), .A(n147), .ZN(n146)
         );
  AOI22_X1 U159 ( .A1(A[1]), .A2(n14), .B1(A[0]), .B2(n20), .ZN(n147) );
  AND3_X1 U160 ( .A1(n97), .A2(n24), .A3(n148), .ZN(n102) );
  MUX2_X1 U161 ( .A(n135), .B(n149), .S(n10), .Z(n144) );
  NOR2_X1 U162 ( .A1(SH[4]), .A2(n150), .ZN(n97) );
  OAI221_X1 U163 ( .B1(n17), .B2(n55), .C1(n105), .C2(n56), .A(n151), .ZN(n96)
         );
  AOI22_X1 U164 ( .A1(A[13]), .A2(n13), .B1(A[12]), .B2(n20), .ZN(n151) );
  NOR2_X1 U165 ( .A1(n24), .A2(n148), .ZN(n114) );
  OAI221_X1 U166 ( .B1(n104), .B2(n59), .C1(n16), .C2(n60), .A(n152), .ZN(n98)
         );
  AOI22_X1 U167 ( .A1(A[9]), .A2(n107), .B1(A[8]), .B2(n20), .ZN(n152) );
  NOR2_X1 U168 ( .A1(n148), .A2(SH[2]), .ZN(n112) );
  OAI221_X1 U169 ( .B1(n18), .B2(n63), .C1(n15), .C2(n64), .A(n153), .ZN(n99)
         );
  AOI22_X1 U170 ( .A1(A[5]), .A2(n14), .B1(A[4]), .B2(n20), .ZN(n153) );
  OR2_X1 U171 ( .A1(n11), .A2(n73), .ZN(n135) );
  MUX2_X1 U172 ( .A(n25), .B(n26), .S(n24), .Z(n73) );
  OAI221_X1 U173 ( .B1(n17), .B2(n51), .C1(n16), .C2(n52), .A(n154), .ZN(n95)
         );
  AOI22_X1 U174 ( .A1(A[17]), .A2(n13), .B1(A[16]), .B2(n20), .ZN(n154) );
  OAI221_X1 U175 ( .B1(n47), .B2(n17), .C1(n15), .C2(n48), .A(n155), .ZN(n94)
         );
  AOI22_X1 U176 ( .A1(A[21]), .A2(n107), .B1(A[20]), .B2(n19), .ZN(n155) );
  NOR2_X1 U177 ( .A1(SH[0]), .A2(SH[1]), .ZN(n108) );
  NOR2_X1 U178 ( .A1(n46), .A2(SH[1]), .ZN(n107) );
  NAND2_X1 U179 ( .A1(n46), .A2(SH[1]), .ZN(n105) );
  NAND2_X1 U180 ( .A1(SH[0]), .A2(SH[1]), .ZN(n104) );
  OR2_X1 U181 ( .A1(SH[6]), .A2(SH[5]), .ZN(n150) );
endmodule


module fpAdder_DW01_sub_3 ( A, B, CI, DIFF, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28;
  wire   [7:1] carry;

  FA_X1 U2_7 ( .A(A[7]), .B(n21), .CI(carry[7]), .S(DIFF[7]) );
  FA_X1 U2_4 ( .A(A[4]), .B(n24), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  FA_X1 U2_0 ( .A(1'b1), .B(A[0]), .CI(n28), .CO(carry[1]), .S(DIFF[0]) );
  XNOR2_X1 U1 ( .A(carry[6]), .B(n1), .ZN(DIFF[6]) );
  XNOR2_X1 U2 ( .A(n22), .B(A[6]), .ZN(n1) );
  NAND2_X1 U3 ( .A1(carry[6]), .A2(n22), .ZN(n2) );
  NAND2_X1 U4 ( .A1(carry[6]), .A2(A[6]), .ZN(n3) );
  NAND2_X1 U5 ( .A1(n22), .A2(A[6]), .ZN(n4) );
  NAND3_X1 U6 ( .A1(n2), .A2(n3), .A3(n4), .ZN(carry[7]) );
  XOR2_X1 U7 ( .A(n25), .B(A[3]), .Z(n5) );
  XOR2_X1 U8 ( .A(carry[3]), .B(n5), .Z(DIFF[3]) );
  NAND2_X1 U9 ( .A1(carry[3]), .A2(n25), .ZN(n6) );
  NAND2_X1 U10 ( .A1(carry[3]), .A2(A[3]), .ZN(n7) );
  NAND2_X1 U11 ( .A1(n25), .A2(A[3]), .ZN(n8) );
  NAND3_X1 U12 ( .A1(n6), .A2(n7), .A3(n8), .ZN(carry[4]) );
  XOR2_X1 U13 ( .A(n23), .B(A[5]), .Z(n9) );
  XOR2_X1 U14 ( .A(carry[5]), .B(n9), .Z(DIFF[5]) );
  NAND2_X1 U15 ( .A1(carry[5]), .A2(n23), .ZN(n10) );
  NAND2_X1 U16 ( .A1(carry[5]), .A2(A[5]), .ZN(n11) );
  NAND2_X1 U17 ( .A1(n23), .A2(A[5]), .ZN(n12) );
  NAND3_X1 U18 ( .A1(n11), .A2(n10), .A3(n12), .ZN(carry[6]) );
  XOR2_X1 U19 ( .A(n26), .B(A[2]), .Z(n13) );
  XOR2_X1 U20 ( .A(carry[2]), .B(n13), .Z(DIFF[2]) );
  NAND2_X1 U21 ( .A1(carry[2]), .A2(n26), .ZN(n14) );
  NAND2_X1 U22 ( .A1(carry[2]), .A2(A[2]), .ZN(n15) );
  NAND2_X1 U23 ( .A1(n26), .A2(A[2]), .ZN(n16) );
  NAND3_X1 U24 ( .A1(n14), .A2(n15), .A3(n16), .ZN(carry[3]) );
  XOR2_X1 U25 ( .A(n27), .B(A[1]), .Z(n17) );
  XOR2_X1 U26 ( .A(carry[1]), .B(n17), .Z(DIFF[1]) );
  NAND2_X1 U27 ( .A1(carry[1]), .A2(n27), .ZN(n18) );
  NAND2_X1 U28 ( .A1(carry[1]), .A2(A[1]), .ZN(n19) );
  NAND2_X1 U29 ( .A1(n27), .A2(A[1]), .ZN(n20) );
  NAND3_X1 U30 ( .A1(n19), .A2(n18), .A3(n20), .ZN(carry[2]) );
  INV_X1 U31 ( .A(B[7]), .ZN(n21) );
  INV_X1 U32 ( .A(B[6]), .ZN(n22) );
  INV_X1 U33 ( .A(B[5]), .ZN(n23) );
  INV_X1 U34 ( .A(B[4]), .ZN(n24) );
  INV_X1 U35 ( .A(B[3]), .ZN(n25) );
  INV_X1 U36 ( .A(B[2]), .ZN(n26) );
  INV_X1 U37 ( .A(B[1]), .ZN(n27) );
  INV_X1 U38 ( .A(B[0]), .ZN(n28) );
endmodule


module fpAdder_DW_rash_1 ( A, DATA_TC, SH, SH_TC, B );
  input [23:0] A;
  input [7:0] SH;
  output [23:0] B;
  input DATA_TC, SH_TC;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148;

  INV_X1 U3 ( .A(SH[2]), .ZN(n17) );
  NOR2_X1 U4 ( .A1(SH[6]), .A2(n4), .ZN(n1) );
  NOR2_X1 U5 ( .A1(SH[6]), .A2(n4), .ZN(n141) );
  NAND2_X1 U6 ( .A1(n104), .A2(n14), .ZN(n65) );
  INV_X1 U7 ( .A(n126), .ZN(n14) );
  INV_X1 U8 ( .A(n68), .ZN(n13) );
  INV_X1 U9 ( .A(SH[0]), .ZN(n39) );
  INV_X1 U10 ( .A(n73), .ZN(n29) );
  INV_X1 U11 ( .A(n83), .ZN(n32) );
  INV_X1 U12 ( .A(n78), .ZN(n24) );
  INV_X1 U13 ( .A(n69), .ZN(n27) );
  INV_X1 U14 ( .A(n77), .ZN(n26) );
  INV_X1 U15 ( .A(n89), .ZN(n22) );
  INV_X1 U16 ( .A(n82), .ZN(n31) );
  INV_X1 U17 ( .A(n87), .ZN(n18) );
  INV_X1 U18 ( .A(SH[7]), .ZN(n15) );
  INV_X1 U19 ( .A(n106), .ZN(n28) );
  INV_X1 U20 ( .A(n116), .ZN(n23) );
  INV_X1 U21 ( .A(n91), .ZN(n21) );
  INV_X1 U22 ( .A(n84), .ZN(n35) );
  INV_X1 U23 ( .A(n81), .ZN(n33) );
  INV_X1 U24 ( .A(n88), .ZN(n19) );
  INV_X1 U25 ( .A(n71), .ZN(n30) );
  INV_X1 U26 ( .A(n76), .ZN(n25) );
  AOI222_X1 U27 ( .A1(n104), .A2(n79), .B1(n105), .B2(n116), .C1(n107), .C2(
        n77), .ZN(n115) );
  AOI222_X1 U28 ( .A1(n104), .A2(n74), .B1(n105), .B2(n106), .C1(n107), .C2(
        n69), .ZN(n103) );
  INV_X1 U29 ( .A(n98), .ZN(n38) );
  INV_X1 U30 ( .A(n85), .ZN(n34) );
  INV_X1 U31 ( .A(n74), .ZN(n37) );
  INV_X1 U32 ( .A(n92), .ZN(n20) );
  INV_X1 U33 ( .A(n79), .ZN(n36) );
  INV_X1 U34 ( .A(A[23]), .ZN(n40) );
  INV_X1 U35 ( .A(A[2]), .ZN(n61) );
  INV_X1 U36 ( .A(A[22]), .ZN(n41) );
  INV_X1 U37 ( .A(A[21]), .ZN(n42) );
  INV_X1 U38 ( .A(A[20]), .ZN(n43) );
  INV_X1 U39 ( .A(A[19]), .ZN(n44) );
  INV_X1 U40 ( .A(A[18]), .ZN(n45) );
  INV_X1 U41 ( .A(A[11]), .ZN(n52) );
  INV_X1 U42 ( .A(A[10]), .ZN(n53) );
  INV_X1 U43 ( .A(A[12]), .ZN(n51) );
  INV_X1 U44 ( .A(A[16]), .ZN(n47) );
  INV_X1 U45 ( .A(A[14]), .ZN(n49) );
  INV_X1 U46 ( .A(A[6]), .ZN(n57) );
  INV_X1 U47 ( .A(A[15]), .ZN(n48) );
  INV_X1 U48 ( .A(A[7]), .ZN(n56) );
  INV_X1 U49 ( .A(A[8]), .ZN(n55) );
  INV_X1 U50 ( .A(A[3]), .ZN(n60) );
  INV_X1 U51 ( .A(A[4]), .ZN(n59) );
  INV_X1 U52 ( .A(A[17]), .ZN(n46) );
  INV_X1 U53 ( .A(A[13]), .ZN(n50) );
  INV_X1 U54 ( .A(A[5]), .ZN(n58) );
  INV_X1 U55 ( .A(A[9]), .ZN(n54) );
  NOR2_X1 U56 ( .A1(SH[4]), .A2(n143), .ZN(n2) );
  INV_X1 U57 ( .A(n1), .ZN(n3) );
  OR2_X1 U58 ( .A1(SH[5]), .A2(SH[3]), .ZN(n4) );
  NOR2_X2 U59 ( .A1(n16), .A2(n17), .ZN(n104) );
  INV_X1 U60 ( .A(n141), .ZN(n16) );
  BUF_X2 U61 ( .A(n101), .Z(n11) );
  BUF_X2 U62 ( .A(n101), .Z(n12) );
  NAND2_X2 U63 ( .A1(n95), .A2(n15), .ZN(n62) );
  NOR2_X1 U64 ( .A1(n39), .A2(SH[1]), .ZN(n5) );
  NOR2_X1 U65 ( .A1(n39), .A2(SH[1]), .ZN(n6) );
  NAND2_X1 U66 ( .A1(n39), .A2(SH[1]), .ZN(n7) );
  NAND2_X1 U67 ( .A1(n39), .A2(SH[1]), .ZN(n8) );
  NAND2_X1 U68 ( .A1(SH[0]), .A2(SH[1]), .ZN(n9) );
  NAND2_X1 U69 ( .A1(SH[0]), .A2(SH[1]), .ZN(n10) );
  OAI222_X1 U70 ( .A1(n35), .A2(n62), .B1(n63), .B2(n64), .C1(n31), .C2(n65), 
        .ZN(B[9]) );
  OAI222_X1 U71 ( .A1(n21), .A2(n62), .B1(n66), .B2(n64), .C1(n22), .C2(n65), 
        .ZN(B[8]) );
  OAI221_X1 U72 ( .B1(n37), .B2(n62), .C1(n28), .C2(n65), .A(n67), .ZN(B[7])
         );
  AOI222_X1 U73 ( .A1(n68), .A2(n69), .B1(n70), .B2(n71), .C1(n72), .C2(n29), 
        .ZN(n67) );
  OAI221_X1 U74 ( .B1(n36), .B2(n62), .C1(n23), .C2(n65), .A(n75), .ZN(B[6])
         );
  AOI222_X1 U75 ( .A1(n72), .A2(n24), .B1(n70), .B2(n76), .C1(n68), .C2(n77), 
        .ZN(n75) );
  OAI221_X1 U76 ( .B1(n34), .B2(n62), .C1(n35), .C2(n65), .A(n80), .ZN(B[5])
         );
  AOI222_X1 U77 ( .A1(n72), .A2(n32), .B1(n70), .B2(n81), .C1(n68), .C2(n82), 
        .ZN(n80) );
  OAI221_X1 U78 ( .B1(n20), .B2(n62), .C1(n21), .C2(n65), .A(n86), .ZN(B[4])
         );
  AOI222_X1 U79 ( .A1(n72), .A2(n87), .B1(n70), .B2(n88), .C1(n68), .C2(n89), 
        .ZN(n86) );
  NOR2_X1 U80 ( .A1(n64), .A2(n17), .ZN(n70) );
  NOR4_X1 U81 ( .A1(n3), .A2(SH[2]), .A3(n2), .A4(SH[7]), .ZN(n72) );
  AOI21_X1 U82 ( .B1(n93), .B2(n94), .A(SH[7]), .ZN(B[3]) );
  NAND2_X1 U83 ( .A1(n95), .A2(n96), .ZN(n94) );
  OAI221_X1 U84 ( .B1(n97), .B2(n57), .C1(n7), .C2(n58), .A(n99), .ZN(n96) );
  AOI22_X1 U85 ( .A1(A[4]), .A2(n6), .B1(A[3]), .B2(n11), .ZN(n99) );
  MUX2_X1 U86 ( .A(n102), .B(n103), .S(n2), .Z(n93) );
  OAI221_X1 U87 ( .B1(n10), .B2(n53), .C1(n98), .C2(n54), .A(n108), .ZN(n74)
         );
  AOI22_X1 U88 ( .A1(A[8]), .A2(n5), .B1(A[7]), .B2(n11), .ZN(n108) );
  OR2_X1 U89 ( .A1(n3), .A2(n109), .ZN(n102) );
  AOI21_X1 U90 ( .B1(n110), .B2(n111), .A(SH[7]), .ZN(B[2]) );
  NAND2_X1 U91 ( .A1(n95), .A2(n112), .ZN(n111) );
  OAI221_X1 U92 ( .B1(n9), .B2(n58), .C1(n8), .C2(n59), .A(n113), .ZN(n112) );
  AOI22_X1 U93 ( .A1(A[3]), .A2(n100), .B1(A[2]), .B2(n11), .ZN(n113) );
  MUX2_X1 U94 ( .A(n114), .B(n115), .S(n2), .Z(n110) );
  OAI221_X1 U95 ( .B1(n97), .B2(n54), .C1(n7), .C2(n55), .A(n117), .ZN(n79) );
  AOI22_X1 U96 ( .A1(A[7]), .A2(n6), .B1(A[6]), .B2(n11), .ZN(n117) );
  NOR2_X1 U97 ( .A1(n62), .A2(n73), .ZN(B[23]) );
  NOR2_X1 U98 ( .A1(n78), .A2(n62), .ZN(B[22]) );
  NOR2_X1 U99 ( .A1(n83), .A2(n62), .ZN(B[21]) );
  NOR2_X1 U100 ( .A1(n18), .A2(n62), .ZN(B[20]) );
  AOI21_X1 U101 ( .B1(n118), .B2(n119), .A(SH[7]), .ZN(B[1]) );
  NAND2_X1 U102 ( .A1(n95), .A2(n120), .ZN(n119) );
  OAI221_X1 U103 ( .B1(n10), .B2(n59), .C1(n98), .C2(n60), .A(n121), .ZN(n120)
         );
  AOI22_X1 U104 ( .A1(A[2]), .A2(n5), .B1(A[1]), .B2(n11), .ZN(n121) );
  MUX2_X1 U105 ( .A(n122), .B(n123), .S(n2), .Z(n118) );
  AOI222_X1 U106 ( .A1(n104), .A2(n85), .B1(n105), .B2(n84), .C1(n107), .C2(
        n82), .ZN(n123) );
  OAI221_X1 U107 ( .B1(n9), .B2(n51), .C1(n8), .C2(n52), .A(n124), .ZN(n84) );
  AOI22_X1 U108 ( .A1(A[10]), .A2(n100), .B1(A[9]), .B2(n11), .ZN(n124) );
  OAI221_X1 U109 ( .B1(n97), .B2(n55), .C1(n7), .C2(n56), .A(n125), .ZN(n85)
         );
  AOI22_X1 U110 ( .A1(A[6]), .A2(n6), .B1(A[5]), .B2(n11), .ZN(n125) );
  NOR3_X1 U111 ( .A1(n3), .A2(n109), .A3(n126), .ZN(B[19]) );
  NOR2_X1 U112 ( .A1(n126), .A2(n114), .ZN(B[18]) );
  OR2_X1 U113 ( .A1(n3), .A2(n127), .ZN(n114) );
  NOR2_X1 U114 ( .A1(n126), .A2(n122), .ZN(B[17]) );
  OR2_X1 U115 ( .A1(n3), .A2(n63), .ZN(n122) );
  MUX2_X1 U116 ( .A(n83), .B(n33), .S(n17), .Z(n63) );
  NOR2_X1 U117 ( .A1(n126), .A2(n128), .ZN(B[16]) );
  OAI222_X1 U118 ( .A1(n27), .A2(n62), .B1(n73), .B2(n13), .C1(n30), .C2(n65), 
        .ZN(B[15]) );
  OAI222_X1 U119 ( .A1(n26), .A2(n62), .B1(n78), .B2(n13), .C1(n25), .C2(n65), 
        .ZN(B[14]) );
  OAI222_X1 U120 ( .A1(n31), .A2(n62), .B1(n83), .B2(n13), .C1(n33), .C2(n65), 
        .ZN(B[13]) );
  OAI221_X1 U121 ( .B1(n10), .B2(n43), .C1(n98), .C2(n44), .A(n129), .ZN(n81)
         );
  AOI22_X1 U122 ( .A1(A[18]), .A2(n5), .B1(A[17]), .B2(n11), .ZN(n129) );
  AOI222_X1 U123 ( .A1(n5), .A2(A[22]), .B1(n38), .B2(A[23]), .C1(n12), .C2(
        A[21]), .ZN(n83) );
  OAI221_X1 U124 ( .B1(n9), .B2(n47), .C1(n8), .C2(n48), .A(n130), .ZN(n82) );
  AOI22_X1 U125 ( .A1(A[14]), .A2(n100), .B1(A[13]), .B2(n11), .ZN(n130) );
  OAI222_X1 U126 ( .A1(n22), .A2(n62), .B1(n18), .B2(n13), .C1(n19), .C2(n65), 
        .ZN(B[12]) );
  NOR2_X1 U127 ( .A1(n64), .A2(SH[2]), .ZN(n68) );
  OAI222_X1 U128 ( .A1(n27), .A2(n65), .B1(n28), .B2(n62), .C1(n109), .C2(n64), 
        .ZN(B[11]) );
  MUX2_X1 U129 ( .A(n73), .B(n30), .S(n17), .Z(n109) );
  OAI221_X1 U130 ( .B1(n41), .B2(n97), .C1(n7), .C2(n42), .A(n131), .ZN(n71)
         );
  AOI22_X1 U131 ( .A1(A[20]), .A2(n6), .B1(A[19]), .B2(n11), .ZN(n131) );
  NAND2_X1 U132 ( .A1(n12), .A2(A[23]), .ZN(n73) );
  OAI221_X1 U133 ( .B1(n97), .B2(n49), .C1(n98), .C2(n50), .A(n132), .ZN(n106)
         );
  AOI22_X1 U134 ( .A1(A[12]), .A2(n5), .B1(A[11]), .B2(n12), .ZN(n132) );
  OAI221_X1 U135 ( .B1(n10), .B2(n45), .C1(n8), .C2(n46), .A(n133), .ZN(n69)
         );
  AOI22_X1 U136 ( .A1(A[16]), .A2(n100), .B1(A[15]), .B2(n12), .ZN(n133) );
  OAI222_X1 U137 ( .A1(n23), .A2(n62), .B1(n127), .B2(n64), .C1(n26), .C2(n65), 
        .ZN(B[10]) );
  OAI221_X1 U138 ( .B1(n9), .B2(n46), .C1(n7), .C2(n47), .A(n134), .ZN(n77) );
  AOI22_X1 U139 ( .A1(A[15]), .A2(n6), .B1(A[14]), .B2(n12), .ZN(n134) );
  NAND2_X1 U140 ( .A1(n14), .A2(n3), .ZN(n64) );
  NAND2_X1 U141 ( .A1(n2), .A2(n15), .ZN(n126) );
  MUX2_X1 U142 ( .A(n78), .B(n25), .S(n17), .Z(n127) );
  OAI221_X1 U143 ( .B1(n42), .B2(n10), .C1(n98), .C2(n43), .A(n135), .ZN(n76)
         );
  AOI22_X1 U144 ( .A1(A[19]), .A2(n5), .B1(A[18]), .B2(n12), .ZN(n135) );
  AOI22_X1 U145 ( .A1(A[22]), .A2(n11), .B1(A[23]), .B2(n6), .ZN(n78) );
  OAI221_X1 U146 ( .B1(n97), .B2(n50), .C1(n8), .C2(n51), .A(n136), .ZN(n116)
         );
  AOI22_X1 U147 ( .A1(A[11]), .A2(n100), .B1(A[10]), .B2(n12), .ZN(n136) );
  AOI21_X1 U148 ( .B1(n137), .B2(n138), .A(SH[7]), .ZN(B[0]) );
  NAND2_X1 U149 ( .A1(n95), .A2(n139), .ZN(n138) );
  OAI221_X1 U150 ( .B1(n10), .B2(n60), .C1(n7), .C2(n61), .A(n140), .ZN(n139)
         );
  AOI22_X1 U151 ( .A1(A[1]), .A2(n6), .B1(A[0]), .B2(n12), .ZN(n140) );
  AND3_X1 U152 ( .A1(n90), .A2(n17), .A3(n1), .ZN(n95) );
  MUX2_X1 U153 ( .A(n128), .B(n142), .S(n2), .Z(n137) );
  NOR2_X1 U154 ( .A1(SH[4]), .A2(n143), .ZN(n90) );
  AOI222_X1 U155 ( .A1(n104), .A2(n92), .B1(n105), .B2(n91), .C1(n107), .C2(
        n89), .ZN(n142) );
  OAI221_X1 U156 ( .B1(n9), .B2(n48), .C1(n98), .C2(n49), .A(n144), .ZN(n89)
         );
  AOI22_X1 U157 ( .A1(A[13]), .A2(n5), .B1(A[12]), .B2(n12), .ZN(n144) );
  NOR2_X1 U158 ( .A1(n17), .A2(n141), .ZN(n107) );
  OAI221_X1 U159 ( .B1(n97), .B2(n52), .C1(n8), .C2(n53), .A(n145), .ZN(n91)
         );
  AOI22_X1 U160 ( .A1(A[9]), .A2(n100), .B1(A[8]), .B2(n12), .ZN(n145) );
  NOR2_X1 U161 ( .A1(SH[2]), .A2(n1), .ZN(n105) );
  OAI221_X1 U162 ( .B1(n10), .B2(n56), .C1(n7), .C2(n57), .A(n146), .ZN(n92)
         );
  AOI22_X1 U163 ( .A1(A[5]), .A2(n6), .B1(A[4]), .B2(n12), .ZN(n146) );
  OR2_X1 U164 ( .A1(n3), .A2(n66), .ZN(n128) );
  MUX2_X1 U165 ( .A(n18), .B(n19), .S(n17), .Z(n66) );
  OAI221_X1 U166 ( .B1(n9), .B2(n44), .C1(n8), .C2(n45), .A(n147), .ZN(n88) );
  AOI22_X1 U167 ( .A1(A[17]), .A2(n5), .B1(A[16]), .B2(n12), .ZN(n147) );
  OAI221_X1 U168 ( .B1(n40), .B2(n9), .C1(n7), .C2(n41), .A(n148), .ZN(n87) );
  AOI22_X1 U169 ( .A1(A[21]), .A2(n100), .B1(A[20]), .B2(n11), .ZN(n148) );
  NOR2_X1 U170 ( .A1(SH[0]), .A2(SH[1]), .ZN(n101) );
  NOR2_X1 U171 ( .A1(n39), .A2(SH[1]), .ZN(n100) );
  NAND2_X1 U172 ( .A1(n39), .A2(SH[1]), .ZN(n98) );
  NAND2_X1 U173 ( .A1(SH[0]), .A2(SH[1]), .ZN(n97) );
  OR2_X1 U174 ( .A1(SH[6]), .A2(SH[5]), .ZN(n143) );
endmodule


module fpAdder_DW01_sub_4 ( A, B, CI, DIFF, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25;
  wire   [7:1] carry;

  FA_X1 U2_7 ( .A(A[7]), .B(n18), .CI(carry[7]), .S(DIFF[7]) );
  FA_X1 U2_5 ( .A(A[5]), .B(n20), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  FA_X1 U2_2 ( .A(A[2]), .B(n23), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  XOR2_X1 U1 ( .A(n22), .B(A[3]), .Z(n1) );
  XOR2_X1 U2 ( .A(n9), .B(n1), .Z(DIFF[3]) );
  NAND2_X1 U3 ( .A1(carry[3]), .A2(n22), .ZN(n2) );
  NAND2_X1 U4 ( .A1(carry[3]), .A2(A[3]), .ZN(n3) );
  NAND2_X1 U5 ( .A1(n22), .A2(A[3]), .ZN(n4) );
  NAND3_X1 U6 ( .A1(n2), .A2(n3), .A3(n4), .ZN(carry[4]) );
  XOR2_X1 U7 ( .A(n21), .B(A[4]), .Z(n5) );
  XOR2_X1 U8 ( .A(carry[4]), .B(n5), .Z(DIFF[4]) );
  NAND2_X1 U9 ( .A1(carry[4]), .A2(n21), .ZN(n6) );
  NAND2_X1 U10 ( .A1(carry[4]), .A2(A[4]), .ZN(n7) );
  NAND2_X1 U11 ( .A1(n21), .A2(A[4]), .ZN(n8) );
  NAND3_X1 U12 ( .A1(n6), .A2(n7), .A3(n8), .ZN(carry[5]) );
  CLKBUF_X1 U13 ( .A(carry[3]), .Z(n9) );
  OR2_X2 U14 ( .A1(n25), .A2(A[0]), .ZN(carry[1]) );
  XOR2_X1 U15 ( .A(n24), .B(A[1]), .Z(n10) );
  XOR2_X1 U16 ( .A(carry[1]), .B(n10), .Z(DIFF[1]) );
  NAND2_X1 U17 ( .A1(carry[1]), .A2(n24), .ZN(n11) );
  NAND2_X1 U18 ( .A1(carry[1]), .A2(A[1]), .ZN(n12) );
  NAND2_X1 U19 ( .A1(n24), .A2(A[1]), .ZN(n13) );
  NAND3_X1 U20 ( .A1(n11), .A2(n12), .A3(n13), .ZN(carry[2]) );
  XNOR2_X1 U21 ( .A(carry[6]), .B(n14), .ZN(DIFF[6]) );
  XNOR2_X1 U22 ( .A(n19), .B(A[6]), .ZN(n14) );
  NAND2_X1 U23 ( .A1(carry[6]), .A2(n19), .ZN(n15) );
  NAND2_X1 U24 ( .A1(carry[6]), .A2(A[6]), .ZN(n16) );
  NAND2_X1 U25 ( .A1(n19), .A2(A[6]), .ZN(n17) );
  NAND3_X1 U26 ( .A1(n15), .A2(n16), .A3(n17), .ZN(carry[7]) );
  XNOR2_X1 U27 ( .A(n25), .B(A[0]), .ZN(DIFF[0]) );
  INV_X1 U28 ( .A(B[7]), .ZN(n18) );
  INV_X1 U29 ( .A(B[6]), .ZN(n19) );
  INV_X1 U30 ( .A(B[5]), .ZN(n20) );
  INV_X1 U31 ( .A(B[4]), .ZN(n21) );
  INV_X1 U32 ( .A(B[3]), .ZN(n22) );
  INV_X1 U33 ( .A(B[2]), .ZN(n23) );
  INV_X1 U34 ( .A(B[1]), .ZN(n24) );
  INV_X1 U35 ( .A(B[0]), .ZN(n25) );
endmodule


module fpAdder_DW01_sub_5 ( A, B, CI, DIFF, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  wire   [7:1] carry;

  FA_X1 U2_5 ( .A(A[5]), .B(n21), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  FA_X1 U2_4 ( .A(A[4]), .B(n22), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  FA_X1 U2_2 ( .A(A[2]), .B(n24), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  INV_X1 U1 ( .A(A[1]), .ZN(n2) );
  XNOR2_X1 U2 ( .A(carry[7]), .B(n1), .ZN(DIFF[7]) );
  XNOR2_X1 U3 ( .A(n21), .B(A[7]), .ZN(n1) );
  OR2_X1 U4 ( .A1(carry[6]), .A2(n5), .ZN(n4) );
  OR2_X1 U5 ( .A1(B[1]), .A2(n2), .ZN(n10) );
  NAND2_X1 U6 ( .A1(carry[6]), .A2(n5), .ZN(n3) );
  NAND2_X1 U7 ( .A1(n3), .A2(n4), .ZN(DIFF[6]) );
  XNOR2_X1 U8 ( .A(n21), .B(A[6]), .ZN(n5) );
  CLKBUF_X1 U9 ( .A(carry[1]), .Z(n6) );
  CLKBUF_X1 U10 ( .A(B[0]), .Z(n7) );
  XOR2_X1 U11 ( .A(n6), .B(A[1]), .Z(n8) );
  XOR2_X1 U12 ( .A(n25), .B(n8), .Z(DIFF[1]) );
  NAND2_X1 U13 ( .A1(n25), .A2(carry[1]), .ZN(n9) );
  NAND2_X1 U14 ( .A1(carry[1]), .A2(A[1]), .ZN(n11) );
  NAND3_X1 U15 ( .A1(n9), .A2(n11), .A3(n10), .ZN(carry[2]) );
  CLKBUF_X1 U16 ( .A(carry[3]), .Z(n12) );
  XOR2_X1 U17 ( .A(n23), .B(A[3]), .Z(n13) );
  XOR2_X1 U18 ( .A(n12), .B(n13), .Z(DIFF[3]) );
  NAND2_X1 U19 ( .A1(carry[3]), .A2(n23), .ZN(n14) );
  NAND2_X1 U20 ( .A1(carry[3]), .A2(A[3]), .ZN(n15) );
  NAND2_X1 U21 ( .A1(n23), .A2(A[3]), .ZN(n16) );
  NAND3_X1 U22 ( .A1(n15), .A2(n14), .A3(n16), .ZN(carry[4]) );
  NAND2_X1 U23 ( .A1(carry[6]), .A2(n21), .ZN(n17) );
  NAND2_X1 U24 ( .A1(carry[6]), .A2(A[6]), .ZN(n18) );
  NAND2_X1 U25 ( .A1(n21), .A2(A[6]), .ZN(n19) );
  NAND3_X1 U26 ( .A1(n18), .A2(n17), .A3(n19), .ZN(carry[7]) );
  XNOR2_X1 U27 ( .A(n26), .B(A[0]), .ZN(DIFF[0]) );
  INV_X1 U28 ( .A(B[4]), .ZN(n22) );
  INV_X1 U29 ( .A(B[3]), .ZN(n23) );
  INV_X1 U30 ( .A(B[2]), .ZN(n24) );
  NAND2_X1 U31 ( .A1(B[0]), .A2(n20), .ZN(carry[1]) );
  INV_X1 U32 ( .A(A[0]), .ZN(n20) );
  INV_X1 U33 ( .A(B[5]), .ZN(n21) );
  INV_X1 U34 ( .A(B[1]), .ZN(n25) );
  INV_X1 U35 ( .A(n7), .ZN(n26) );
endmodule


module fpAdder ( clk, reset, enable, A, B, result, overFlow );
  input [31:0] A;
  input [31:0] B;
  output [31:0] result;
  input clk, reset, enable;
  output overFlow;
  wire   IBA, IBB, N135, N137, N138, N139, N140, N141, N142, N143, N144, N145,
         N146, N147, N148, N149, N150, N151, N152, N153, N154, N155, N156,
         N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167,
         N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178,
         N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189,
         N190, N191, N192, N193, N194, N195, N196, N197, N198, N199, N200,
         N201, N202, N203, N204, N205, N206, N207, N208, N212, N213, N214,
         N215, N216, N217, N218, N219, N220, N221, N222, N223, N224, N225,
         N226, N227, N228, N229, N230, N231, N232, N233, N234, N235, N236,
         N238, N239, N240, N241, N242, N243, N244, N245, N278, N280, N281,
         N282, N283, N284, N285, N286, N287, N288, N289, N290, N291, N292,
         N293, N294, N295, N296, N297, N298, N299, N300, N301, N302, N303,
         N304, N305, N306, N307, N308, N309, N310, N311, N312, N313, N314,
         N315, N316, N317, N318, N319, N320, N321, N322, N323, N324, N325,
         N326, N327, N480, N481, N482, N483, N484, N518, N519, N521, N549,
         N550, N551, N552, N553, N554, N555, N556, N557, N558, N559, N560,
         N561, N562, N563, N564, N565, N566, N567, N568, N569, N570, N571,
         N580, N581, N582, N583, N584, N585, N586, N587, N612, n74, n76, n1350,
         n136, n1370, n1380, n1390, n1400, n1410, n1420, n1430, n1440, n1450,
         n1460, n1470, n1480, n1490, n1500, n1510, n1520, n1530, n1540, n1550,
         n1560, n1570, n1580, n1590, n1600, n1610, n1620, n1630, n1640, n1650,
         n1660, n1670, n1680, n1690, n1700, n1710, n1720, n1730, n1740, n1750,
         n1760, n1770, n1780, n1790, n1800, n1810, n1820, n1830, n1840, n1850,
         n1860, n1870, n1880, n1890, n1900, n1910, n1920, n1930, n1940, n1950,
         n1960, n1980, n1990, n2000, n2010, n2020, n2030, n2040, n2050, n2060,
         n2070, n209, n210, n211, n2120, n2130, n2140, n2150, n2160, n2170,
         n2180, n2190, n2200, n2210, n2220, n2230, n2240, n2250, n2260, n2270,
         n2280, n2290, n2300, n2310, n2320, n2330, n2340, n2350, n2360, n237,
         n2380, n2390, n2400, n2410, n2420, n2430, n2440, n2450, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n2780, n279, n2800, n2810,
         n2820, n2830, n2840, n2850, n2860, n2870, n2880, n2890, n2900, n2910,
         n2920, n2930, n2940, n2950, n2960, n2970, n2980, n2990, n3000, n3010,
         n3020, n3030, n3040, n3050, n3060, n3070, n3080, n3090, n3100, n3110,
         n3120, n3130, n3140, n3150, n3160, n3170, n3180, n3190, n3200, n3210,
         n3220, n3230, n3240, n3250, n3260, n3270, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n4800, n4810, n4820, n4830, n4840, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, N576, N575,
         r145_B_23_, sll_78_ML_int_5__16_, sll_78_ML_int_5__17_,
         sll_78_ML_int_5__18_, sll_78_ML_int_5__19_, sll_78_ML_int_5__20_,
         sll_78_ML_int_5__21_, sll_78_ML_int_5__22_, sll_78_ML_int_4__8_,
         sll_78_ML_int_4__9_, sll_78_ML_int_4__10_, sll_78_ML_int_4__11_,
         sll_78_ML_int_4__12_, sll_78_ML_int_4__13_, sll_78_ML_int_4__14_,
         sll_78_ML_int_4__15_, sll_78_ML_int_4__16_, sll_78_ML_int_4__17_,
         sll_78_ML_int_4__18_, sll_78_ML_int_4__19_, sll_78_ML_int_4__20_,
         sll_78_ML_int_4__21_, sll_78_ML_int_4__22_, sll_78_ML_int_3__0_,
         sll_78_ML_int_3__1_, sll_78_ML_int_3__2_, sll_78_ML_int_3__3_,
         sll_78_ML_int_3__4_, sll_78_ML_int_3__5_, sll_78_ML_int_3__6_,
         sll_78_ML_int_3__7_, sll_78_ML_int_3__8_, sll_78_ML_int_3__9_,
         sll_78_ML_int_3__10_, sll_78_ML_int_3__11_, sll_78_ML_int_3__12_,
         sll_78_ML_int_3__13_, sll_78_ML_int_3__14_, sll_78_ML_int_3__15_,
         sll_78_ML_int_3__16_, sll_78_ML_int_3__17_, sll_78_ML_int_3__18_,
         sll_78_ML_int_3__19_, sll_78_ML_int_3__20_, sll_78_ML_int_3__21_,
         sll_78_ML_int_3__22_, sll_78_ML_int_2__0_, sll_78_ML_int_2__1_,
         sll_78_ML_int_2__2_, sll_78_ML_int_2__3_, sll_78_ML_int_2__4_,
         sll_78_ML_int_2__5_, sll_78_ML_int_2__6_, sll_78_ML_int_2__7_,
         sll_78_ML_int_2__8_, sll_78_ML_int_2__9_, sll_78_ML_int_2__10_,
         sll_78_ML_int_2__11_, sll_78_ML_int_2__12_, sll_78_ML_int_2__13_,
         sll_78_ML_int_2__14_, sll_78_ML_int_2__15_, sll_78_ML_int_2__16_,
         sll_78_ML_int_2__17_, sll_78_ML_int_2__18_, sll_78_ML_int_2__19_,
         sll_78_ML_int_2__20_, sll_78_ML_int_2__21_, sll_78_ML_int_2__22_,
         sll_78_ML_int_1__0_, sll_78_ML_int_1__1_, sll_78_ML_int_1__2_,
         sll_78_ML_int_1__3_, sll_78_ML_int_1__4_, sll_78_ML_int_1__5_,
         sll_78_ML_int_1__6_, sll_78_ML_int_1__7_, sll_78_ML_int_1__8_,
         sll_78_ML_int_1__9_, sll_78_ML_int_1__10_, sll_78_ML_int_1__11_,
         sll_78_ML_int_1__12_, sll_78_ML_int_1__13_, sll_78_ML_int_1__14_,
         sll_78_ML_int_1__15_, sll_78_ML_int_1__16_, sll_78_ML_int_1__17_,
         sll_78_ML_int_1__18_, sll_78_ML_int_1__19_, sll_78_ML_int_1__20_,
         sll_78_ML_int_1__21_, sll_78_ML_int_1__22_, sll_78_A_0_, sll_78_A_1_,
         sll_78_A_2_, sll_78_A_3_, sll_78_A_4_, sll_78_A_5_, sll_78_A_6_,
         sll_78_A_7_, sll_78_A_8_, sll_78_A_9_, sll_78_A_10_, sll_78_A_11_,
         sll_78_A_12_, sll_78_A_13_, sll_78_A_14_, sll_78_A_15_, sll_78_A_16_,
         sll_78_A_17_, sll_78_A_18_, sll_78_A_19_, sll_78_A_20_, sll_78_A_21_,
         sll_78_A_22_, sub_78_B_1_, sub_78_B_2_, sub_78_B_4_, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n5180, n5190,
         n520, n5210, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n5490, n5500, n5510, n5520,
         n5530, n5540, n5550, n5560, n5570, n5580, n5590, n5600, n5610, n5620,
         n5630, n5640, n5650, n5660, n5670, n5680, n5690, n5700, n5710, n572,
         n573, n574, n5750, n5760, n577, n578, n579, n5800, n5810, n5820,
         n5830, n5840, n5850, n5860, n5870, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n6120, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766;
  wire   [30:0] A_reg;
  wire   [31:0] B_reg;
  wire   [23:0] MB;
  wire   [22:0] MA;
  wire   [4:0] MSB;

  DFF_X1 B_reg_reg_31_ ( .D(n505), .CK(clk), .Q(B_reg[31]), .QN(n74) );
  DFF_X1 B_reg_reg_30_ ( .D(n504), .CK(clk), .Q(B_reg[30]), .QN(n76) );
  DFF_X1 B_reg_reg_29_ ( .D(n503), .CK(clk), .Q(B_reg[29]), .QN(n1350) );
  DFF_X1 B_reg_reg_28_ ( .D(n502), .CK(clk), .Q(B_reg[28]), .QN(n136) );
  DFF_X1 B_reg_reg_27_ ( .D(n501), .CK(clk), .Q(B_reg[27]), .QN(n1370) );
  DFF_X1 B_reg_reg_25_ ( .D(n499), .CK(clk), .Q(B_reg[25]), .QN(n1390) );
  DFF_X1 B_reg_reg_24_ ( .D(n498), .CK(clk), .Q(B_reg[24]), .QN(n1400) );
  DFF_X1 B_reg_reg_23_ ( .D(n497), .CK(clk), .Q(B_reg[23]), .QN(n1410) );
  DFF_X1 B_reg_reg_22_ ( .D(n496), .CK(clk), .Q(B_reg[22]), .QN(n1420) );
  DFF_X1 B_reg_reg_21_ ( .D(n495), .CK(clk), .Q(B_reg[21]), .QN(n1430) );
  DFF_X1 B_reg_reg_20_ ( .D(n494), .CK(clk), .Q(B_reg[20]), .QN(n1440) );
  DFF_X1 B_reg_reg_19_ ( .D(n493), .CK(clk), .Q(B_reg[19]), .QN(n1450) );
  DFF_X1 B_reg_reg_18_ ( .D(n492), .CK(clk), .Q(B_reg[18]), .QN(n1460) );
  DFF_X1 B_reg_reg_17_ ( .D(n491), .CK(clk), .Q(B_reg[17]), .QN(n1470) );
  DFF_X1 B_reg_reg_16_ ( .D(n490), .CK(clk), .Q(B_reg[16]), .QN(n1480) );
  DFF_X1 B_reg_reg_15_ ( .D(n489), .CK(clk), .Q(B_reg[15]), .QN(n1490) );
  DFF_X1 B_reg_reg_14_ ( .D(n488), .CK(clk), .Q(B_reg[14]), .QN(n1500) );
  DFF_X1 B_reg_reg_13_ ( .D(n487), .CK(clk), .Q(B_reg[13]), .QN(n1510) );
  DFF_X1 B_reg_reg_12_ ( .D(n486), .CK(clk), .Q(B_reg[12]), .QN(n1520) );
  DFF_X1 B_reg_reg_11_ ( .D(n485), .CK(clk), .Q(B_reg[11]), .QN(n1530) );
  DFF_X1 B_reg_reg_10_ ( .D(n4840), .CK(clk), .Q(B_reg[10]), .QN(n1540) );
  DFF_X1 B_reg_reg_9_ ( .D(n4830), .CK(clk), .Q(B_reg[9]), .QN(n1550) );
  DFF_X1 B_reg_reg_8_ ( .D(n4820), .CK(clk), .Q(B_reg[8]), .QN(n1560) );
  DFF_X1 B_reg_reg_7_ ( .D(n4810), .CK(clk), .Q(B_reg[7]), .QN(n1570) );
  DFF_X1 B_reg_reg_6_ ( .D(n4800), .CK(clk), .Q(B_reg[6]), .QN(n1580) );
  DFF_X1 B_reg_reg_5_ ( .D(n479), .CK(clk), .Q(B_reg[5]), .QN(n1590) );
  DFF_X1 B_reg_reg_4_ ( .D(n478), .CK(clk), .Q(B_reg[4]), .QN(n1600) );
  DFF_X1 B_reg_reg_3_ ( .D(n477), .CK(clk), .Q(B_reg[3]), .QN(n1610) );
  DFF_X1 B_reg_reg_2_ ( .D(n476), .CK(clk), .Q(B_reg[2]), .QN(n1620) );
  DFF_X1 B_reg_reg_1_ ( .D(n475), .CK(clk), .Q(B_reg[1]), .QN(n1630) );
  DFF_X1 B_reg_reg_0_ ( .D(n474), .CK(clk), .Q(B_reg[0]), .QN(n1640) );
  DFF_X1 A_reg_reg_31_ ( .D(n473), .CK(clk), .QN(n1650) );
  DFF_X1 A_reg_reg_30_ ( .D(n472), .CK(clk), .Q(A_reg[30]), .QN(n1660) );
  DFF_X1 A_reg_reg_29_ ( .D(n471), .CK(clk), .Q(A_reg[29]), .QN(n1670) );
  DFF_X1 A_reg_reg_28_ ( .D(n470), .CK(clk), .Q(A_reg[28]), .QN(n1680) );
  DFF_X1 A_reg_reg_27_ ( .D(n469), .CK(clk), .Q(A_reg[27]), .QN(n1690) );
  DFF_X1 A_reg_reg_26_ ( .D(n468), .CK(clk), .Q(A_reg[26]), .QN(n1700) );
  DFF_X1 A_reg_reg_25_ ( .D(n467), .CK(clk), .Q(A_reg[25]), .QN(n1710) );
  DFF_X1 A_reg_reg_24_ ( .D(n466), .CK(clk), .Q(A_reg[24]), .QN(n1720) );
  DFF_X1 A_reg_reg_23_ ( .D(n465), .CK(clk), .Q(A_reg[23]), .QN(n1730) );
  DFF_X1 A_reg_reg_22_ ( .D(n464), .CK(clk), .Q(A_reg[22]), .QN(n1740) );
  DFF_X1 A_reg_reg_21_ ( .D(n463), .CK(clk), .Q(A_reg[21]), .QN(n1750) );
  DFF_X1 A_reg_reg_20_ ( .D(n462), .CK(clk), .Q(A_reg[20]), .QN(n1760) );
  DFF_X1 A_reg_reg_19_ ( .D(n461), .CK(clk), .Q(A_reg[19]), .QN(n1770) );
  DFF_X1 A_reg_reg_18_ ( .D(n460), .CK(clk), .Q(A_reg[18]), .QN(n1780) );
  DFF_X1 A_reg_reg_17_ ( .D(n459), .CK(clk), .Q(A_reg[17]), .QN(n1790) );
  DFF_X1 A_reg_reg_16_ ( .D(n458), .CK(clk), .Q(A_reg[16]), .QN(n1800) );
  DFF_X1 A_reg_reg_15_ ( .D(n457), .CK(clk), .Q(A_reg[15]), .QN(n1810) );
  DFF_X1 A_reg_reg_14_ ( .D(n456), .CK(clk), .Q(A_reg[14]), .QN(n1820) );
  DFF_X1 A_reg_reg_13_ ( .D(n455), .CK(clk), .Q(A_reg[13]), .QN(n1830) );
  DFF_X1 A_reg_reg_12_ ( .D(n454), .CK(clk), .Q(A_reg[12]), .QN(n1840) );
  DFF_X1 A_reg_reg_11_ ( .D(n453), .CK(clk), .Q(A_reg[11]), .QN(n1850) );
  DFF_X1 A_reg_reg_10_ ( .D(n452), .CK(clk), .Q(A_reg[10]), .QN(n1860) );
  DFF_X1 A_reg_reg_9_ ( .D(n451), .CK(clk), .Q(A_reg[9]), .QN(n1870) );
  DFF_X1 A_reg_reg_8_ ( .D(n450), .CK(clk), .Q(A_reg[8]), .QN(n1880) );
  DFF_X1 A_reg_reg_7_ ( .D(n449), .CK(clk), .Q(A_reg[7]), .QN(n1890) );
  DFF_X1 A_reg_reg_6_ ( .D(n448), .CK(clk), .Q(A_reg[6]), .QN(n1900) );
  DFF_X1 A_reg_reg_5_ ( .D(n447), .CK(clk), .Q(A_reg[5]), .QN(n1910) );
  DFF_X1 A_reg_reg_4_ ( .D(n446), .CK(clk), .Q(A_reg[4]), .QN(n1920) );
  DFF_X1 A_reg_reg_3_ ( .D(n445), .CK(clk), .Q(A_reg[3]), .QN(n1930) );
  DFF_X1 A_reg_reg_2_ ( .D(n444), .CK(clk), .Q(A_reg[2]), .QN(n1940) );
  DFF_X1 A_reg_reg_1_ ( .D(n443), .CK(clk), .Q(A_reg[1]), .QN(n1950) );
  DFF_X1 A_reg_reg_0_ ( .D(n442), .CK(clk), .Q(A_reg[0]), .QN(n1960) );
  DLH_X1 MSB_reg_4_ ( .G(N612), .D(N484), .Q(MSB[4]) );
  DLH_X1 MSB_reg_3_ ( .G(N612), .D(N483), .Q(MSB[3]) );
  DLH_X1 MSB_reg_2_ ( .G(N612), .D(N482), .Q(MSB[2]) );
  DLH_X1 MSB_reg_1_ ( .G(N612), .D(N481), .Q(MSB[1]) );
  DLH_X1 MSB_reg_0_ ( .G(N612), .D(N480), .Q(MSB[0]) );
  AND2_X2 U95 ( .A1(n529), .A2(N236), .ZN(n2070) );
  OAI21_X2 U359 ( .B1(n5800), .B2(n1630), .A(n415), .ZN(MB[1]) );
  fpAdder_DW01_sub_1 sub_70 ( .A(MB), .B({r145_B_23_, MA}), .CI(1'b0), .DIFF({
        N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, 
        N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304}) );
  fpAdder_DW01_sub_2 sub_68 ( .A({r145_B_23_, MA[22:1], n528}), .B(MB), .CI(
        1'b0), .DIFF({N303, N302, N301, N300, N299, N298, N297, N296, N295, 
        N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, 
        N282, N281, N280}) );
  fpAdder_DW01_inc_0 add_63 ( .A({N208, N207, N206, N205, N204, N203, N202, 
        N201}), .SUM({N245, N244, N243, N242, N241, N240, N239, N238}) );
  fpAdder_DW01_add_0 add_59 ( .A({1'b0, r145_B_23_, MA[22:1], n528}), .B({1'b0, 
        MB[23:1], n5180}), .CI(1'b0), .SUM({N236, N235, N234, N233, N232, N231, 
        N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, 
        N218, N217, N216, N215, N214, N213, N212}) );
  fpAdder_DW_rash_0 srl_52 ( .A({IBB, B_reg[22:0]}), .DATA_TC(1'b0), .SH({N144, 
        N143, N142, N141, N140, N139, N138, N137}), .SH_TC(1'b0), .B({N168, 
        N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, 
        N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145}) );
  fpAdder_DW01_sub_3 sub_52 ( .A(A_reg[30:23]), .B(B_reg[30:23]), .CI(1'b0), 
        .DIFF({N144, N143, N142, N141, N140, N139, N138, N137}) );
  fpAdder_DW_rash_1 srl_55 ( .A({IBA, A_reg[22:0]}), .DATA_TC(1'b0), .SH({N176, 
        N175, N174, N173, N172, N171, N170, N169}), .SH_TC(1'b0), .B({N200, 
        N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, 
        N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177}) );
  fpAdder_DW01_sub_4 sub_55 ( .A({B_reg[30:24], n531}), .B(A_reg[30:23]), .CI(
        1'b0), .DIFF({N176, N175, N174, N173, N172, N171, N170, N169}) );
  fpAdder_DW01_sub_5 sub_79_2 ( .A({N208, N207, N206, N205, N204, N203, N202, 
        N201}), .B({n5190, n5190, n5190, N576, n525, n345, n344, n527}), .CI(
        1'b0), .DIFF({N587, N586, N585, N584, N583, N582, N581, N580}) );
  MUX2_X1 sll_78_M1_0_1 ( .A(sll_78_A_1_), .B(sll_78_A_0_), .S(n510), .Z(
        sll_78_ML_int_1__1_) );
  MUX2_X1 sll_78_M1_0_2 ( .A(sll_78_A_2_), .B(sll_78_A_1_), .S(n510), .Z(
        sll_78_ML_int_1__2_) );
  MUX2_X1 sll_78_M1_0_3 ( .A(sll_78_A_3_), .B(sll_78_A_2_), .S(n510), .Z(
        sll_78_ML_int_1__3_) );
  MUX2_X1 sll_78_M1_0_4 ( .A(sll_78_A_4_), .B(sll_78_A_3_), .S(n510), .Z(
        sll_78_ML_int_1__4_) );
  MUX2_X1 sll_78_M1_0_5 ( .A(sll_78_A_5_), .B(sll_78_A_4_), .S(n510), .Z(
        sll_78_ML_int_1__5_) );
  MUX2_X1 sll_78_M1_0_6 ( .A(sll_78_A_6_), .B(sll_78_A_5_), .S(n510), .Z(
        sll_78_ML_int_1__6_) );
  MUX2_X1 sll_78_M1_0_7 ( .A(sll_78_A_7_), .B(sll_78_A_6_), .S(n510), .Z(
        sll_78_ML_int_1__7_) );
  MUX2_X1 sll_78_M1_0_8 ( .A(sll_78_A_8_), .B(sll_78_A_7_), .S(n510), .Z(
        sll_78_ML_int_1__8_) );
  MUX2_X1 sll_78_M1_0_9 ( .A(sll_78_A_9_), .B(sll_78_A_8_), .S(n510), .Z(
        sll_78_ML_int_1__9_) );
  MUX2_X1 sll_78_M1_0_10 ( .A(sll_78_A_10_), .B(sll_78_A_9_), .S(n510), .Z(
        sll_78_ML_int_1__10_) );
  MUX2_X1 sll_78_M1_0_11 ( .A(sll_78_A_11_), .B(sll_78_A_10_), .S(n510), .Z(
        sll_78_ML_int_1__11_) );
  MUX2_X1 sll_78_M1_0_12 ( .A(sll_78_A_12_), .B(sll_78_A_11_), .S(n510), .Z(
        sll_78_ML_int_1__12_) );
  MUX2_X1 sll_78_M1_0_13 ( .A(sll_78_A_13_), .B(sll_78_A_12_), .S(n510), .Z(
        sll_78_ML_int_1__13_) );
  MUX2_X1 sll_78_M1_0_14 ( .A(sll_78_A_14_), .B(sll_78_A_13_), .S(n510), .Z(
        sll_78_ML_int_1__14_) );
  MUX2_X1 sll_78_M1_0_15 ( .A(sll_78_A_15_), .B(sll_78_A_14_), .S(n510), .Z(
        sll_78_ML_int_1__15_) );
  MUX2_X1 sll_78_M1_0_16 ( .A(sll_78_A_16_), .B(sll_78_A_15_), .S(n510), .Z(
        sll_78_ML_int_1__16_) );
  MUX2_X1 sll_78_M1_0_17 ( .A(sll_78_A_17_), .B(sll_78_A_16_), .S(n510), .Z(
        sll_78_ML_int_1__17_) );
  MUX2_X1 sll_78_M1_0_18 ( .A(sll_78_A_18_), .B(sll_78_A_17_), .S(n510), .Z(
        sll_78_ML_int_1__18_) );
  MUX2_X1 sll_78_M1_0_19 ( .A(sll_78_A_19_), .B(sll_78_A_18_), .S(n510), .Z(
        sll_78_ML_int_1__19_) );
  MUX2_X1 sll_78_M1_0_20 ( .A(sll_78_A_20_), .B(sll_78_A_19_), .S(n510), .Z(
        sll_78_ML_int_1__20_) );
  MUX2_X1 sll_78_M1_0_21 ( .A(sll_78_A_21_), .B(sll_78_A_20_), .S(n510), .Z(
        sll_78_ML_int_1__21_) );
  MUX2_X1 sll_78_M1_0_22 ( .A(sll_78_A_22_), .B(sll_78_A_21_), .S(n510), .Z(
        sll_78_ML_int_1__22_) );
  MUX2_X1 sll_78_M1_1_2 ( .A(sll_78_ML_int_1__2_), .B(sll_78_ML_int_1__0_), 
        .S(N518), .Z(sll_78_ML_int_2__2_) );
  MUX2_X1 sll_78_M1_1_3 ( .A(sll_78_ML_int_1__3_), .B(sll_78_ML_int_1__1_), 
        .S(N518), .Z(sll_78_ML_int_2__3_) );
  MUX2_X1 sll_78_M1_1_4 ( .A(sll_78_ML_int_1__4_), .B(sll_78_ML_int_1__2_), 
        .S(N518), .Z(sll_78_ML_int_2__4_) );
  MUX2_X1 sll_78_M1_1_5 ( .A(sll_78_ML_int_1__5_), .B(sll_78_ML_int_1__3_), 
        .S(N518), .Z(sll_78_ML_int_2__5_) );
  MUX2_X1 sll_78_M1_1_6 ( .A(sll_78_ML_int_1__6_), .B(sll_78_ML_int_1__4_), 
        .S(N518), .Z(sll_78_ML_int_2__6_) );
  MUX2_X1 sll_78_M1_1_7 ( .A(sll_78_ML_int_1__7_), .B(sll_78_ML_int_1__5_), 
        .S(N518), .Z(sll_78_ML_int_2__7_) );
  MUX2_X1 sll_78_M1_1_8 ( .A(sll_78_ML_int_1__8_), .B(sll_78_ML_int_1__6_), 
        .S(N518), .Z(sll_78_ML_int_2__8_) );
  MUX2_X1 sll_78_M1_1_9 ( .A(sll_78_ML_int_1__9_), .B(sll_78_ML_int_1__7_), 
        .S(N518), .Z(sll_78_ML_int_2__9_) );
  MUX2_X1 sll_78_M1_1_10 ( .A(sll_78_ML_int_1__10_), .B(sll_78_ML_int_1__8_), 
        .S(N518), .Z(sll_78_ML_int_2__10_) );
  MUX2_X1 sll_78_M1_1_11 ( .A(sll_78_ML_int_1__11_), .B(sll_78_ML_int_1__9_), 
        .S(N518), .Z(sll_78_ML_int_2__11_) );
  MUX2_X1 sll_78_M1_1_12 ( .A(sll_78_ML_int_1__12_), .B(sll_78_ML_int_1__10_), 
        .S(N518), .Z(sll_78_ML_int_2__12_) );
  MUX2_X1 sll_78_M1_1_13 ( .A(sll_78_ML_int_1__13_), .B(sll_78_ML_int_1__11_), 
        .S(N518), .Z(sll_78_ML_int_2__13_) );
  MUX2_X1 sll_78_M1_1_14 ( .A(sll_78_ML_int_1__14_), .B(sll_78_ML_int_1__12_), 
        .S(N518), .Z(sll_78_ML_int_2__14_) );
  MUX2_X1 sll_78_M1_1_15 ( .A(sll_78_ML_int_1__15_), .B(sll_78_ML_int_1__13_), 
        .S(N518), .Z(sll_78_ML_int_2__15_) );
  MUX2_X1 sll_78_M1_1_16 ( .A(sll_78_ML_int_1__16_), .B(sll_78_ML_int_1__14_), 
        .S(N518), .Z(sll_78_ML_int_2__16_) );
  MUX2_X1 sll_78_M1_1_17 ( .A(sll_78_ML_int_1__17_), .B(sll_78_ML_int_1__15_), 
        .S(N518), .Z(sll_78_ML_int_2__17_) );
  MUX2_X1 sll_78_M1_1_18 ( .A(sll_78_ML_int_1__18_), .B(sll_78_ML_int_1__16_), 
        .S(N518), .Z(sll_78_ML_int_2__18_) );
  MUX2_X1 sll_78_M1_1_19 ( .A(sll_78_ML_int_1__19_), .B(sll_78_ML_int_1__17_), 
        .S(N518), .Z(sll_78_ML_int_2__19_) );
  MUX2_X1 sll_78_M1_1_20 ( .A(sll_78_ML_int_1__20_), .B(sll_78_ML_int_1__18_), 
        .S(N518), .Z(sll_78_ML_int_2__20_) );
  MUX2_X1 sll_78_M1_1_21 ( .A(sll_78_ML_int_1__21_), .B(sll_78_ML_int_1__19_), 
        .S(N518), .Z(sll_78_ML_int_2__21_) );
  MUX2_X1 sll_78_M1_1_22 ( .A(sll_78_ML_int_1__22_), .B(sll_78_ML_int_1__20_), 
        .S(N518), .Z(sll_78_ML_int_2__22_) );
  MUX2_X1 sll_78_M1_2_4 ( .A(sll_78_ML_int_2__4_), .B(sll_78_ML_int_2__0_), 
        .S(N519), .Z(sll_78_ML_int_3__4_) );
  MUX2_X1 sll_78_M1_2_5 ( .A(sll_78_ML_int_2__5_), .B(sll_78_ML_int_2__1_), 
        .S(N519), .Z(sll_78_ML_int_3__5_) );
  MUX2_X1 sll_78_M1_2_6 ( .A(sll_78_ML_int_2__6_), .B(sll_78_ML_int_2__2_), 
        .S(N519), .Z(sll_78_ML_int_3__6_) );
  MUX2_X1 sll_78_M1_2_7 ( .A(sll_78_ML_int_2__7_), .B(sll_78_ML_int_2__3_), 
        .S(N519), .Z(sll_78_ML_int_3__7_) );
  MUX2_X1 sll_78_M1_2_8 ( .A(sll_78_ML_int_2__8_), .B(sll_78_ML_int_2__4_), 
        .S(N519), .Z(sll_78_ML_int_3__8_) );
  MUX2_X1 sll_78_M1_2_9 ( .A(sll_78_ML_int_2__9_), .B(sll_78_ML_int_2__5_), 
        .S(N519), .Z(sll_78_ML_int_3__9_) );
  MUX2_X1 sll_78_M1_2_10 ( .A(sll_78_ML_int_2__10_), .B(sll_78_ML_int_2__6_), 
        .S(N519), .Z(sll_78_ML_int_3__10_) );
  MUX2_X1 sll_78_M1_2_11 ( .A(sll_78_ML_int_2__11_), .B(sll_78_ML_int_2__7_), 
        .S(N519), .Z(sll_78_ML_int_3__11_) );
  MUX2_X1 sll_78_M1_2_12 ( .A(sll_78_ML_int_2__12_), .B(sll_78_ML_int_2__8_), 
        .S(N519), .Z(sll_78_ML_int_3__12_) );
  MUX2_X1 sll_78_M1_2_13 ( .A(sll_78_ML_int_2__13_), .B(sll_78_ML_int_2__9_), 
        .S(N519), .Z(sll_78_ML_int_3__13_) );
  MUX2_X1 sll_78_M1_2_14 ( .A(sll_78_ML_int_2__14_), .B(sll_78_ML_int_2__10_), 
        .S(N519), .Z(sll_78_ML_int_3__14_) );
  MUX2_X1 sll_78_M1_2_15 ( .A(sll_78_ML_int_2__15_), .B(sll_78_ML_int_2__11_), 
        .S(N519), .Z(sll_78_ML_int_3__15_) );
  MUX2_X1 sll_78_M1_2_16 ( .A(sll_78_ML_int_2__16_), .B(sll_78_ML_int_2__12_), 
        .S(N519), .Z(sll_78_ML_int_3__16_) );
  MUX2_X1 sll_78_M1_2_17 ( .A(sll_78_ML_int_2__17_), .B(sll_78_ML_int_2__13_), 
        .S(N519), .Z(sll_78_ML_int_3__17_) );
  MUX2_X1 sll_78_M1_2_18 ( .A(sll_78_ML_int_2__18_), .B(sll_78_ML_int_2__14_), 
        .S(N519), .Z(sll_78_ML_int_3__18_) );
  MUX2_X1 sll_78_M1_2_19 ( .A(sll_78_ML_int_2__19_), .B(sll_78_ML_int_2__15_), 
        .S(N519), .Z(sll_78_ML_int_3__19_) );
  MUX2_X1 sll_78_M1_2_20 ( .A(sll_78_ML_int_2__20_), .B(sll_78_ML_int_2__16_), 
        .S(N519), .Z(sll_78_ML_int_3__20_) );
  MUX2_X1 sll_78_M1_2_21 ( .A(sll_78_ML_int_2__21_), .B(sll_78_ML_int_2__17_), 
        .S(N519), .Z(sll_78_ML_int_3__21_) );
  MUX2_X1 sll_78_M1_2_22 ( .A(sll_78_ML_int_2__22_), .B(sll_78_ML_int_2__18_), 
        .S(N519), .Z(sll_78_ML_int_3__22_) );
  MUX2_X1 sll_78_M1_3_8 ( .A(sll_78_ML_int_3__8_), .B(sll_78_ML_int_3__0_), 
        .S(n526), .Z(sll_78_ML_int_4__8_) );
  MUX2_X1 sll_78_M1_3_9 ( .A(sll_78_ML_int_3__9_), .B(sll_78_ML_int_3__1_), 
        .S(n526), .Z(sll_78_ML_int_4__9_) );
  MUX2_X1 sll_78_M1_3_10 ( .A(sll_78_ML_int_3__10_), .B(sll_78_ML_int_3__2_), 
        .S(n526), .Z(sll_78_ML_int_4__10_) );
  MUX2_X1 sll_78_M1_3_11 ( .A(sll_78_ML_int_3__11_), .B(sll_78_ML_int_3__3_), 
        .S(n526), .Z(sll_78_ML_int_4__11_) );
  MUX2_X1 sll_78_M1_3_12 ( .A(sll_78_ML_int_3__12_), .B(sll_78_ML_int_3__4_), 
        .S(N575), .Z(sll_78_ML_int_4__12_) );
  MUX2_X1 sll_78_M1_3_13 ( .A(sll_78_ML_int_3__13_), .B(sll_78_ML_int_3__5_), 
        .S(n526), .Z(sll_78_ML_int_4__13_) );
  MUX2_X1 sll_78_M1_3_14 ( .A(sll_78_ML_int_3__14_), .B(sll_78_ML_int_3__6_), 
        .S(N575), .Z(sll_78_ML_int_4__14_) );
  MUX2_X1 sll_78_M1_3_15 ( .A(sll_78_ML_int_3__15_), .B(sll_78_ML_int_3__7_), 
        .S(N575), .Z(sll_78_ML_int_4__15_) );
  MUX2_X1 sll_78_M1_3_16 ( .A(sll_78_ML_int_3__16_), .B(sll_78_ML_int_3__8_), 
        .S(N575), .Z(sll_78_ML_int_4__16_) );
  MUX2_X1 sll_78_M1_3_17 ( .A(sll_78_ML_int_3__17_), .B(sll_78_ML_int_3__9_), 
        .S(n526), .Z(sll_78_ML_int_4__17_) );
  MUX2_X1 sll_78_M1_3_18 ( .A(sll_78_ML_int_3__18_), .B(sll_78_ML_int_3__10_), 
        .S(n526), .Z(sll_78_ML_int_4__18_) );
  MUX2_X1 sll_78_M1_3_19 ( .A(sll_78_ML_int_3__19_), .B(sll_78_ML_int_3__11_), 
        .S(n526), .Z(sll_78_ML_int_4__19_) );
  MUX2_X1 sll_78_M1_3_20 ( .A(sll_78_ML_int_3__20_), .B(sll_78_ML_int_3__12_), 
        .S(n526), .Z(sll_78_ML_int_4__20_) );
  MUX2_X1 sll_78_M1_3_21 ( .A(sll_78_ML_int_3__21_), .B(sll_78_ML_int_3__13_), 
        .S(n526), .Z(sll_78_ML_int_4__21_) );
  MUX2_X1 sll_78_M1_3_22 ( .A(sll_78_ML_int_3__22_), .B(sll_78_ML_int_3__14_), 
        .S(n526), .Z(sll_78_ML_int_4__22_) );
  MUX2_X1 sll_78_M1_4_16 ( .A(sll_78_ML_int_4__16_), .B(n614), .S(N521), .Z(
        sll_78_ML_int_5__16_) );
  MUX2_X1 sll_78_M1_4_17 ( .A(sll_78_ML_int_4__17_), .B(n610), .S(N521), .Z(
        sll_78_ML_int_5__17_) );
  MUX2_X1 sll_78_M1_4_18 ( .A(sll_78_ML_int_4__18_), .B(n6120), .S(N521), .Z(
        sll_78_ML_int_5__18_) );
  MUX2_X1 sll_78_M1_4_19 ( .A(sll_78_ML_int_4__19_), .B(n608), .S(N521), .Z(
        sll_78_ML_int_5__19_) );
  MUX2_X1 sll_78_M1_4_20 ( .A(sll_78_ML_int_4__20_), .B(n613), .S(N521), .Z(
        sll_78_ML_int_5__20_) );
  MUX2_X1 sll_78_M1_4_21 ( .A(sll_78_ML_int_4__21_), .B(n609), .S(N521), .Z(
        sll_78_ML_int_5__21_) );
  MUX2_X1 sll_78_M1_4_22 ( .A(sll_78_ML_int_4__22_), .B(n611), .S(N521), .Z(
        sll_78_ML_int_5__22_) );
  DFF_X1 result_reg_31_ ( .D(n738), .CK(clk), .Q(result[31]) );
  DFF_X1 result_reg_23_ ( .D(n439), .CK(clk), .Q(result[23]) );
  DFF_X1 result_reg_24_ ( .D(n438), .CK(clk), .Q(result[24]) );
  DFF_X1 result_reg_25_ ( .D(n437), .CK(clk), .Q(result[25]) );
  DFF_X1 result_reg_26_ ( .D(n436), .CK(clk), .Q(result[26]) );
  DFF_X1 result_reg_27_ ( .D(n435), .CK(clk), .Q(result[27]) );
  DFF_X1 result_reg_28_ ( .D(n434), .CK(clk), .Q(result[28]) );
  DFF_X1 result_reg_29_ ( .D(n433), .CK(clk), .Q(result[29]) );
  DFF_X1 result_reg_30_ ( .D(n432), .CK(clk), .Q(result[30]) );
  DFF_X1 overFlow_reg ( .D(n441), .CK(clk), .Q(overFlow) );
  DFF_X1 result_reg_0_ ( .D(n440), .CK(clk), .Q(result[0]) );
  DFF_X1 result_reg_21_ ( .D(n523), .CK(clk), .Q(result[21]) );
  DFF_X1 result_reg_2_ ( .D(n524), .CK(clk), .Q(result[2]) );
  DFF_X1 result_reg_18_ ( .D(n729), .CK(clk), .Q(result[18]) );
  DFF_X1 result_reg_17_ ( .D(n727), .CK(clk), .Q(result[17]) );
  DFF_X1 result_reg_6_ ( .D(n705), .CK(clk), .Q(result[6]) );
  DFF_X1 result_reg_19_ ( .D(n731), .CK(clk), .Q(result[19]) );
  DFF_X1 result_reg_16_ ( .D(n725), .CK(clk), .Q(result[16]) );
  DFF_X1 result_reg_13_ ( .D(n719), .CK(clk), .Q(result[13]) );
  DFF_X1 result_reg_10_ ( .D(n713), .CK(clk), .Q(result[10]) );
  DFF_X1 result_reg_7_ ( .D(n707), .CK(clk), .Q(result[7]) );
  DFF_X1 result_reg_4_ ( .D(n701), .CK(clk), .Q(result[4]) );
  DFF_X1 result_reg_1_ ( .D(n696), .CK(clk), .Q(result[1]) );
  DFF_X1 result_reg_15_ ( .D(n723), .CK(clk), .Q(result[15]) );
  DFF_X1 result_reg_14_ ( .D(n721), .CK(clk), .Q(result[14]) );
  DFF_X1 result_reg_3_ ( .D(n699), .CK(clk), .Q(result[3]) );
  DFF_X1 result_reg_22_ ( .D(n736), .CK(clk), .Q(result[22]) );
  DFF_X1 result_reg_20_ ( .D(n733), .CK(clk), .Q(result[20]) );
  DFF_X1 result_reg_12_ ( .D(n717), .CK(clk), .Q(result[12]) );
  DFF_X1 result_reg_11_ ( .D(n715), .CK(clk), .Q(result[11]) );
  DFF_X1 result_reg_8_ ( .D(n709), .CK(clk), .Q(result[8]) );
  DFF_X1 result_reg_5_ ( .D(n703), .CK(clk), .Q(result[5]) );
  DFF_X1 result_reg_9_ ( .D(n711), .CK(clk), .Q(result[9]) );
  DFF_X1 B_reg_reg_26_ ( .D(n500), .CK(clk), .Q(B_reg[26]), .QN(n1380) );
  NAND2_X1 U518 ( .A1(n380), .A2(n379), .ZN(n506) );
  NAND3_X1 U519 ( .A1(n381), .A2(n378), .A3(n507), .ZN(n358) );
  INV_X1 U520 ( .A(n506), .ZN(n507) );
  OR2_X2 U521 ( .A1(n511), .A2(n262), .ZN(n513) );
  OAI21_X2 U522 ( .B1(n579), .B2(n1640), .A(n426), .ZN(MB[0]) );
  BUF_X1 U523 ( .A(n594), .Z(n593) );
  BUF_X1 U524 ( .A(n594), .Z(n592) );
  INV_X1 U525 ( .A(n592), .ZN(n5750) );
  INV_X1 U526 ( .A(n593), .ZN(n579) );
  OAI21_X1 U527 ( .B1(n5800), .B2(n1490), .A(n420), .ZN(MB[15]) );
  AOI22_X1 U528 ( .A1(N309), .A2(n5700), .B1(N285), .B2(N278), .ZN(n375) );
  OAI22_X1 U529 ( .A1(n578), .A2(n757), .B1(n5840), .B2(n1880), .ZN(MA[8]) );
  OAI21_X1 U530 ( .B1(n579), .B2(n1560), .A(n404), .ZN(MB[8]) );
  OAI22_X1 U531 ( .A1(n577), .A2(n749), .B1(n591), .B2(n1850), .ZN(MA[11]) );
  OAI22_X1 U532 ( .A1(n577), .A2(n750), .B1(n591), .B2(n1840), .ZN(MA[12]) );
  OAI21_X1 U533 ( .B1(n5810), .B2(n1520), .A(n423), .ZN(MB[12]) );
  OAI22_X1 U534 ( .A1(n577), .A2(n754), .B1(n588), .B2(n1760), .ZN(MA[20]) );
  OAI22_X1 U535 ( .A1(n578), .A2(n745), .B1(n5860), .B2(n1930), .ZN(MA[3]) );
  OAI21_X1 U536 ( .B1(n579), .B2(n1610), .A(n409), .ZN(MB[3]) );
  OAI22_X1 U537 ( .A1(n577), .A2(n752), .B1(n590), .B2(n1820), .ZN(MA[14]) );
  OAI22_X1 U538 ( .A1(n578), .A2(n753), .B1(n590), .B2(n1810), .ZN(MA[15]) );
  OAI21_X1 U539 ( .B1(n5810), .B2(n1540), .A(n425), .ZN(MB[10]) );
  OAI21_X1 U540 ( .B1(n579), .B2(n1580), .A(n406), .ZN(MB[6]) );
  OAI22_X1 U541 ( .A1(n577), .A2(n760), .B1(n589), .B2(n1790), .ZN(MA[17]) );
  OAI21_X1 U542 ( .B1(n5800), .B2(n1470), .A(n418), .ZN(MB[17]) );
  OAI22_X1 U543 ( .A1(n577), .A2(n761), .B1(n589), .B2(n1780), .ZN(MA[18]) );
  OAI21_X1 U544 ( .B1(n5800), .B2(n1460), .A(n417), .ZN(MB[18]) );
  OAI22_X1 U545 ( .A1(n578), .A2(n1350), .B1(n5830), .B2(n1670), .ZN(N207) );
  OAI22_X1 U546 ( .A1(n578), .A2(n1380), .B1(n5840), .B2(n1700), .ZN(N204) );
  OAI22_X1 U547 ( .A1(n577), .A2(n756), .B1(n5870), .B2(n1740), .ZN(MA[22]) );
  OAI21_X1 U548 ( .B1(n5800), .B2(n1430), .A(n413), .ZN(MB[21]) );
  OAI21_X1 U549 ( .B1(n5800), .B2(n1440), .A(n414), .ZN(MB[20]) );
  AOI22_X1 U550 ( .A1(N319), .A2(n5660), .B1(N295), .B2(n5630), .ZN(n371) );
  XNOR2_X1 U551 ( .A(n1650), .B(B_reg[31]), .ZN(n254) );
  AOI22_X1 U552 ( .A1(N323), .A2(n5650), .B1(N299), .B2(n5630), .ZN(n355) );
  INV_X1 U553 ( .A(n514), .ZN(N484) );
  NAND2_X1 U554 ( .A1(sub_78_B_4_), .A2(n526), .ZN(n508) );
  BUF_X1 U555 ( .A(n573), .Z(n572) );
  INV_X1 U556 ( .A(n343), .ZN(n509) );
  INV_X2 U557 ( .A(n509), .ZN(n510) );
  OR2_X1 U558 ( .A1(n2010), .A2(n1980), .ZN(n511) );
  NOR2_X1 U559 ( .A1(n261), .A2(n513), .ZN(n512) );
  AND2_X2 U560 ( .A1(n517), .A2(n740), .ZN(n543) );
  AND2_X2 U561 ( .A1(n517), .A2(n740), .ZN(n2050) );
  OAI22_X4 U562 ( .A1(n578), .A2(n1400), .B1(n1720), .B2(n5820), .ZN(N202) );
  OAI21_X1 U563 ( .B1(n5800), .B2(n1620), .A(n410), .ZN(MB[2]) );
  AOI21_X1 U564 ( .B1(n342), .B2(MSB[0]), .A(N480), .ZN(n343) );
  AND4_X2 U565 ( .A1(n357), .A2(n355), .A3(n356), .A4(n354), .ZN(n514) );
  CLKBUF_X1 U566 ( .A(n1410), .Z(n515) );
  AND2_X2 U567 ( .A1(n517), .A2(n740), .ZN(n544) );
  AND2_X1 U568 ( .A1(n259), .A2(n512), .ZN(n516) );
  AND2_X1 U569 ( .A1(n260), .A2(n259), .ZN(n255) );
  BUF_X2 U570 ( .A(MA[0]), .Z(n528) );
  OAI22_X2 U571 ( .A1(n578), .A2(n747), .B1(n588), .B2(n1950), .ZN(MA[1]) );
  BUF_X1 U572 ( .A(n529), .Z(n517) );
  CLKBUF_X1 U573 ( .A(MB[0]), .Z(n5180) );
  NOR2_X1 U574 ( .A1(n261), .A2(n513), .ZN(n260) );
  INV_X2 U575 ( .A(n593), .ZN(n577) );
  CLKBUF_X1 U576 ( .A(n573), .Z(n5700) );
  CLKBUF_X1 U577 ( .A(n573), .Z(n5710) );
  CLKBUF_X1 U578 ( .A(n595), .Z(n5870) );
  AND2_X1 U579 ( .A1(sub_78_B_4_), .A2(N575), .ZN(n5190) );
  CLKBUF_X1 U580 ( .A(n378), .Z(n520) );
  AND2_X1 U581 ( .A1(n252), .A2(N236), .ZN(n5210) );
  AND2_X1 U582 ( .A1(n252), .A2(N236), .ZN(n522) );
  INV_X1 U583 ( .A(n572), .ZN(n5630) );
  INV_X1 U584 ( .A(n592), .ZN(n5760) );
  INV_X1 U585 ( .A(n593), .ZN(n578) );
  INV_X1 U586 ( .A(n593), .ZN(n5800) );
  NOR3_X1 U587 ( .A1(sll_78_A_17_), .A2(sll_78_A_19_), .A3(sll_78_A_18_), .ZN(
        n367) );
  INV_X1 U588 ( .A(n604), .ZN(n607) );
  BUF_X1 U589 ( .A(n573), .Z(n5660) );
  BUF_X1 U590 ( .A(n573), .Z(n5650) );
  BUF_X1 U591 ( .A(n5650), .Z(n5670) );
  BUF_X1 U592 ( .A(n5640), .Z(n5690) );
  BUF_X1 U593 ( .A(n5660), .Z(n5680) );
  NOR2_X1 U594 ( .A1(sll_78_A_7_), .A2(sll_78_A_6_), .ZN(n389) );
  BUF_X1 U595 ( .A(n573), .Z(n5640) );
  INV_X1 U596 ( .A(n602), .ZN(n609) );
  INV_X1 U597 ( .A(N521), .ZN(n606) );
  AOI21_X1 U598 ( .B1(n394), .B2(n379), .A(sll_78_A_21_), .ZN(n393) );
  OAI21_X1 U599 ( .B1(sll_78_A_18_), .B2(n395), .A(n355), .ZN(n394) );
  AOI21_X1 U600 ( .B1(n396), .B2(n366), .A(sll_78_A_17_), .ZN(n395) );
  NAND4_X1 U601 ( .A1(n368), .A2(n369), .A3(n370), .A4(n371), .ZN(n363) );
  NAND4_X1 U602 ( .A1(n374), .A2(n375), .A3(n376), .A4(n377), .ZN(n353) );
  NOR3_X1 U603 ( .A1(n351), .A2(n352), .A3(n353), .ZN(n350) );
  AOI211_X1 U604 ( .C1(n384), .C2(n385), .A(sll_78_A_19_), .B(sll_78_A_18_), 
        .ZN(n382) );
  NAND2_X1 U605 ( .A1(n379), .A2(n380), .ZN(n383) );
  NOR2_X1 U606 ( .A1(sll_78_A_17_), .A2(sll_78_A_16_), .ZN(n384) );
  NAND4_X1 U607 ( .A1(n359), .A2(n360), .A3(n361), .A4(n362), .ZN(n351) );
  NOR2_X1 U608 ( .A1(sll_78_A_8_), .A2(n363), .ZN(n362) );
  OAI211_X1 U609 ( .C1(n386), .C2(n387), .A(n370), .B(n371), .ZN(n385) );
  NAND2_X1 U610 ( .A1(n368), .A2(n369), .ZN(n387) );
  NOR3_X1 U611 ( .A1(n388), .A2(sll_78_A_11_), .A3(sll_78_A_10_), .ZN(n386) );
  AOI211_X1 U612 ( .C1(n389), .C2(n390), .A(sll_78_A_9_), .B(sll_78_A_8_), 
        .ZN(n388) );
  NAND3_X1 U613 ( .A1(n374), .A2(n375), .A3(n352), .ZN(n390) );
  INV_X1 U614 ( .A(n359), .ZN(sll_78_A_10_) );
  INV_X1 U615 ( .A(n354), .ZN(sll_78_A_18_) );
  INV_X1 U616 ( .A(n361), .ZN(sll_78_A_9_) );
  INV_X1 U617 ( .A(n356), .ZN(sll_78_A_17_) );
  OAI21_X1 U618 ( .B1(sll_78_A_6_), .B2(n401), .A(n377), .ZN(n400) );
  AOI21_X1 U619 ( .B1(n402), .B2(n374), .A(sll_78_A_5_), .ZN(n401) );
  OAI21_X1 U620 ( .B1(sll_78_A_2_), .B2(n348), .A(n392), .ZN(n402) );
  OAI21_X1 U621 ( .B1(sll_78_A_14_), .B2(n397), .A(n371), .ZN(n396) );
  AOI21_X1 U622 ( .B1(n398), .B2(n368), .A(sll_78_A_13_), .ZN(n397) );
  OAI21_X1 U623 ( .B1(sll_78_A_10_), .B2(n399), .A(n360), .ZN(n398) );
  AOI21_X1 U624 ( .B1(n400), .B2(n373), .A(sll_78_A_9_), .ZN(n399) );
  NAND2_X1 U625 ( .A1(n391), .A2(n392), .ZN(n352) );
  INV_X1 U626 ( .A(n360), .ZN(sll_78_A_11_) );
  BUF_X1 U627 ( .A(n595), .Z(n588) );
  BUF_X1 U628 ( .A(n596), .Z(n5860) );
  BUF_X1 U629 ( .A(n596), .Z(n5840) );
  BUF_X1 U630 ( .A(n595), .Z(n591) );
  BUF_X1 U631 ( .A(n595), .Z(n590) );
  CLKBUF_X1 U632 ( .A(n590), .Z(n589) );
  INV_X1 U633 ( .A(N278), .ZN(n573) );
  INV_X1 U634 ( .A(n373), .ZN(sll_78_A_8_) );
  INV_X1 U635 ( .A(N236), .ZN(n740) );
  INV_X1 U636 ( .A(n355), .ZN(sll_78_A_19_) );
  INV_X1 U637 ( .A(n376), .ZN(sll_78_A_6_) );
  BUF_X1 U638 ( .A(n596), .Z(n5850) );
  INV_X1 U639 ( .A(n366), .ZN(sll_78_A_16_) );
  INV_X1 U640 ( .A(n377), .ZN(sll_78_A_7_) );
  INV_X1 U641 ( .A(n370), .ZN(sll_78_A_14_) );
  INV_X1 U642 ( .A(n369), .ZN(sll_78_A_13_) );
  INV_X1 U643 ( .A(n375), .ZN(sll_78_A_5_) );
  NAND2_X1 U644 ( .A1(n353), .A2(n373), .ZN(n372) );
  INV_X1 U645 ( .A(n380), .ZN(sll_78_A_21_) );
  INV_X1 U646 ( .A(n371), .ZN(sll_78_A_15_) );
  INV_X1 U647 ( .A(n368), .ZN(sll_78_A_12_) );
  INV_X1 U648 ( .A(n374), .ZN(sll_78_A_4_) );
  INV_X1 U649 ( .A(n391), .ZN(sll_78_A_2_) );
  INV_X1 U650 ( .A(n379), .ZN(sll_78_A_20_) );
  INV_X1 U651 ( .A(n392), .ZN(sll_78_A_3_) );
  NAND2_X1 U652 ( .A1(n739), .A2(n364), .ZN(N482) );
  OAI211_X1 U653 ( .C1(n365), .C2(n363), .A(n366), .B(n367), .ZN(n364) );
  NOR4_X1 U654 ( .A1(n372), .A2(sll_78_A_9_), .A3(sll_78_A_11_), .A4(
        sll_78_A_10_), .ZN(n365) );
  INV_X1 U655 ( .A(n348), .ZN(sll_78_A_1_) );
  INV_X1 U656 ( .A(n381), .ZN(sll_78_A_22_) );
  INV_X1 U657 ( .A(n349), .ZN(sll_78_A_0_) );
  BUF_X1 U658 ( .A(n589), .Z(n5820) );
  BUF_X1 U659 ( .A(n589), .Z(n5830) );
  INV_X1 U660 ( .A(MB[23]), .ZN(n655) );
  INV_X1 U661 ( .A(n648), .ZN(n695) );
  XNOR2_X1 U662 ( .A(n347), .B(n605), .ZN(N521) );
  AOI22_X1 U663 ( .A1(N316), .A2(n5670), .B1(N292), .B2(n5630), .ZN(n368) );
  AOI22_X1 U664 ( .A1(N308), .A2(n5700), .B1(N284), .B2(N278), .ZN(n374) );
  AOI22_X1 U665 ( .A1(N324), .A2(n5650), .B1(N300), .B2(n5630), .ZN(n379) );
  AOI22_X1 U666 ( .A1(N311), .A2(n5690), .B1(N287), .B2(N278), .ZN(n377) );
  AOI22_X1 U667 ( .A1(N318), .A2(n5660), .B1(N294), .B2(n5630), .ZN(n370) );
  AOI22_X1 U668 ( .A1(N312), .A2(n5690), .B1(N288), .B2(N278), .ZN(n373) );
  AOI22_X1 U669 ( .A1(N320), .A2(n5660), .B1(N296), .B2(n5630), .ZN(n366) );
  AOI22_X1 U670 ( .A1(N317), .A2(n5670), .B1(N293), .B2(n5630), .ZN(n369) );
  AOI22_X1 U671 ( .A1(N307), .A2(n5700), .B1(N283), .B2(n5630), .ZN(n392) );
  AOI22_X1 U672 ( .A1(N315), .A2(n5670), .B1(N291), .B2(N278), .ZN(n360) );
  AOI22_X1 U673 ( .A1(N325), .A2(n5640), .B1(N301), .B2(n5630), .ZN(n380) );
  AOI22_X1 U674 ( .A1(N305), .A2(n5710), .B1(N281), .B2(N278), .ZN(n348) );
  AOI22_X1 U675 ( .A1(N326), .A2(n5640), .B1(N302), .B2(n5630), .ZN(n381) );
  AOI22_X1 U676 ( .A1(N313), .A2(n5680), .B1(N289), .B2(N278), .ZN(n361) );
  AOI22_X1 U677 ( .A1(N310), .A2(n5690), .B1(N286), .B2(N278), .ZN(n376) );
  AOI22_X1 U678 ( .A1(N306), .A2(n5710), .B1(N282), .B2(n5630), .ZN(n391) );
  AOI22_X1 U679 ( .A1(N314), .A2(n5680), .B1(N290), .B2(N278), .ZN(n359) );
  AOI22_X1 U680 ( .A1(N304), .A2(n5710), .B1(N280), .B2(N278), .ZN(n349) );
  AOI22_X1 U681 ( .A1(N321), .A2(n5650), .B1(N297), .B2(n5630), .ZN(n356) );
  AOI22_X1 U682 ( .A1(N322), .A2(n5680), .B1(N298), .B2(n5630), .ZN(n354) );
  BUF_X1 U683 ( .A(n2040), .Z(n542) );
  BUF_X2 U684 ( .A(n2040), .Z(n540) );
  BUF_X2 U685 ( .A(n2040), .Z(n541) );
  INV_X1 U686 ( .A(n600), .ZN(n608) );
  INV_X1 U687 ( .A(n599), .ZN(n6120) );
  INV_X1 U688 ( .A(n598), .ZN(n610) );
  INV_X1 U689 ( .A(n603), .ZN(n611) );
  INV_X1 U690 ( .A(n597), .ZN(n614) );
  INV_X1 U691 ( .A(n601), .ZN(n613) );
  BUF_X1 U692 ( .A(n545), .Z(n547) );
  BUF_X1 U693 ( .A(n545), .Z(n548) );
  BUF_X1 U694 ( .A(n545), .Z(n5490) );
  BUF_X1 U695 ( .A(n546), .Z(n5500) );
  BUF_X1 U696 ( .A(n546), .Z(n5510) );
  BUF_X1 U697 ( .A(n5530), .Z(n5570) );
  BUF_X1 U698 ( .A(n5540), .Z(n5580) );
  BUF_X1 U699 ( .A(n5540), .Z(n5590) );
  BUF_X1 U700 ( .A(n5530), .Z(n5560) );
  BUF_X1 U701 ( .A(n5530), .Z(n5550) );
  NOR2_X1 U702 ( .A1(n740), .A2(n254), .ZN(n258) );
  NOR2_X1 U703 ( .A1(n254), .A2(N236), .ZN(n263) );
  AOI222_X1 U704 ( .A1(N582), .A2(n254), .B1(n263), .B2(N203), .C1(N240), .C2(
        n258), .ZN(n267) );
  AOI222_X1 U705 ( .A1(N583), .A2(n254), .B1(n263), .B2(N204), .C1(N241), .C2(
        n258), .ZN(n266) );
  AOI222_X1 U706 ( .A1(N584), .A2(n254), .B1(n263), .B2(N205), .C1(N242), .C2(
        n258), .ZN(n265) );
  AOI222_X1 U707 ( .A1(N585), .A2(n254), .B1(n263), .B2(N206), .C1(N243), .C2(
        n258), .ZN(n264) );
  OAI21_X1 U708 ( .B1(n5800), .B2(n766), .A(n411), .ZN(MB[23]) );
  INV_X1 U709 ( .A(IBB), .ZN(n766) );
  NAND2_X1 U710 ( .A1(N168), .A2(n5760), .ZN(n411) );
  AOI222_X1 U711 ( .A1(N580), .A2(n254), .B1(n263), .B2(N201), .C1(N238), .C2(
        n258), .ZN(n2010) );
  AOI222_X1 U712 ( .A1(N581), .A2(n254), .B1(n263), .B2(N202), .C1(N239), .C2(
        n258), .ZN(n1980) );
  AOI222_X1 U713 ( .A1(N586), .A2(n254), .B1(n263), .B2(N207), .C1(N244), .C2(
        n258), .ZN(n262) );
  INV_X1 U714 ( .A(n646), .ZN(n694) );
  INV_X1 U715 ( .A(MB[22]), .ZN(n656) );
  INV_X1 U716 ( .A(sub_78_B_1_), .ZN(N518) );
  INV_X1 U717 ( .A(sub_78_B_2_), .ZN(N519) );
  INV_X1 U718 ( .A(MA[17]), .ZN(n675) );
  INV_X1 U719 ( .A(MA[16]), .ZN(n676) );
  INV_X1 U720 ( .A(MA[18]), .ZN(n674) );
  INV_X1 U721 ( .A(MA[19]), .ZN(n673) );
  INV_X1 U722 ( .A(MA[21]), .ZN(n679) );
  INV_X1 U723 ( .A(MA[20]), .ZN(n680) );
  INV_X1 U724 ( .A(MA[15]), .ZN(n681) );
  INV_X1 U725 ( .A(MA[14]), .ZN(n682) );
  INV_X1 U726 ( .A(MA[5]), .ZN(n692) );
  INV_X1 U727 ( .A(MA[4]), .ZN(n693) );
  INV_X1 U728 ( .A(MA[3]), .ZN(n689) );
  INV_X1 U729 ( .A(MA[2]), .ZN(n688) );
  INV_X1 U730 ( .A(MA[9]), .ZN(n677) );
  INV_X1 U731 ( .A(MA[8]), .ZN(n678) );
  INV_X1 U732 ( .A(MA[7]), .ZN(n690) );
  INV_X1 U733 ( .A(MA[6]), .ZN(n691) );
  INV_X1 U734 ( .A(MA[13]), .ZN(n683) );
  INV_X1 U735 ( .A(MA[12]), .ZN(n684) );
  INV_X1 U736 ( .A(MA[11]), .ZN(n685) );
  INV_X1 U737 ( .A(MA[10]), .ZN(n686) );
  INV_X1 U738 ( .A(MA[1]), .ZN(n687) );
  INV_X1 U739 ( .A(n427), .ZN(r145_B_23_) );
  AOI22_X1 U740 ( .A1(n5820), .A2(N200), .B1(IBA), .B2(n5750), .ZN(n427) );
  XNOR2_X1 U741 ( .A(n347), .B(n346), .ZN(N576) );
  NOR4_X1 U742 ( .A1(n264), .A2(n265), .A3(n266), .A4(n267), .ZN(n259) );
  INV_X1 U743 ( .A(MB[1]), .ZN(n665) );
  INV_X1 U744 ( .A(MB[10]), .ZN(n664) );
  INV_X1 U745 ( .A(MB[15]), .ZN(n659) );
  INV_X1 U746 ( .A(MB[17]), .ZN(n651) );
  INV_X1 U747 ( .A(MB[19]), .ZN(n649) );
  INV_X1 U748 ( .A(MB[21]), .ZN(n657) );
  INV_X1 U749 ( .A(MB[5]), .ZN(n670) );
  INV_X1 U750 ( .A(MB[7]), .ZN(n668) );
  INV_X1 U751 ( .A(MB[3]), .ZN(n667) );
  INV_X1 U752 ( .A(MB[14]), .ZN(n660) );
  INV_X1 U753 ( .A(MB[4]), .ZN(n671) );
  INV_X1 U754 ( .A(MB[2]), .ZN(n666) );
  INV_X1 U755 ( .A(MB[16]), .ZN(n652) );
  INV_X1 U756 ( .A(MB[18]), .ZN(n650) );
  INV_X1 U757 ( .A(MB[20]), .ZN(n658) );
  INV_X1 U758 ( .A(MB[8]), .ZN(n654) );
  INV_X1 U759 ( .A(MB[6]), .ZN(n669) );
  INV_X1 U760 ( .A(MB[13]), .ZN(n661) );
  INV_X1 U761 ( .A(MB[11]), .ZN(n663) );
  INV_X1 U762 ( .A(MB[12]), .ZN(n662) );
  INV_X1 U763 ( .A(MB[9]), .ZN(n653) );
  OR3_X1 U764 ( .A1(n534), .A2(n535), .A3(n735), .ZN(n523) );
  OR3_X1 U765 ( .A1(n536), .A2(n537), .A3(n698), .ZN(n524) );
  BUF_X1 U766 ( .A(n2000), .Z(n5620) );
  INV_X1 U767 ( .A(n254), .ZN(n765) );
  BUF_X1 U768 ( .A(n2000), .Z(n5610) );
  BUF_X1 U769 ( .A(n2000), .Z(n5600) );
  INV_X1 U770 ( .A(N192), .ZN(n753) );
  OAI22_X1 U771 ( .A1(n577), .A2(n751), .B1(n591), .B2(n1830), .ZN(MA[13]) );
  INV_X1 U772 ( .A(N190), .ZN(n751) );
  INV_X1 U773 ( .A(N188), .ZN(n749) );
  OAI22_X1 U774 ( .A1(n578), .A2(n748), .B1(n592), .B2(n1860), .ZN(MA[10]) );
  INV_X1 U775 ( .A(N187), .ZN(n748) );
  INV_X1 U776 ( .A(N178), .ZN(n747) );
  OAI22_X1 U777 ( .A1(n578), .A2(n742), .B1(n5850), .B2(n1910), .ZN(MA[5]) );
  INV_X1 U778 ( .A(N182), .ZN(n742) );
  INV_X1 U779 ( .A(N180), .ZN(n745) );
  OAI22_X1 U780 ( .A1(n579), .A2(n744), .B1(n5860), .B2(n1890), .ZN(MA[7]) );
  INV_X1 U781 ( .A(N184), .ZN(n744) );
  INV_X1 U782 ( .A(N194), .ZN(n760) );
  OAI22_X1 U783 ( .A1(n577), .A2(n762), .B1(n589), .B2(n1770), .ZN(MA[19]) );
  INV_X1 U784 ( .A(N196), .ZN(n762) );
  OAI22_X1 U785 ( .A1(n578), .A2(n755), .B1(n5870), .B2(n1750), .ZN(MA[21]) );
  INV_X1 U786 ( .A(N198), .ZN(n755) );
  INV_X1 U787 ( .A(N191), .ZN(n752) );
  INV_X1 U788 ( .A(N189), .ZN(n750) );
  OAI22_X1 U789 ( .A1(n578), .A2(n758), .B1(n5840), .B2(n1870), .ZN(MA[9]) );
  INV_X1 U790 ( .A(N186), .ZN(n758) );
  OAI22_X1 U791 ( .A1(n577), .A2(n741), .B1(n5870), .B2(n1920), .ZN(MA[4]) );
  INV_X1 U792 ( .A(N181), .ZN(n741) );
  OAI22_X1 U793 ( .A1(n577), .A2(n743), .B1(n5850), .B2(n1900), .ZN(MA[6]) );
  INV_X1 U794 ( .A(N183), .ZN(n743) );
  INV_X1 U795 ( .A(N185), .ZN(n757) );
  OAI22_X1 U796 ( .A1(n579), .A2(n759), .B1(n590), .B2(n1800), .ZN(MA[16]) );
  INV_X1 U797 ( .A(N193), .ZN(n759) );
  INV_X1 U798 ( .A(N195), .ZN(n761) );
  INV_X1 U799 ( .A(N197), .ZN(n754) );
  INV_X1 U800 ( .A(N199), .ZN(n756) );
  OAI21_X1 U801 ( .B1(n5800), .B2(n1500), .A(n421), .ZN(MB[14]) );
  NAND2_X1 U802 ( .A1(N159), .A2(n5750), .ZN(n421) );
  OAI21_X1 U803 ( .B1(n5800), .B2(n1480), .A(n419), .ZN(MB[16]) );
  NAND2_X1 U804 ( .A1(N161), .A2(n5760), .ZN(n419) );
  NAND2_X1 U805 ( .A1(N163), .A2(n5760), .ZN(n417) );
  NAND2_X1 U806 ( .A1(N165), .A2(n5760), .ZN(n414) );
  NAND2_X1 U807 ( .A1(N153), .A2(n5750), .ZN(n404) );
  NAND2_X1 U808 ( .A1(N146), .A2(n5750), .ZN(n415) );
  NAND2_X1 U809 ( .A1(N157), .A2(n5760), .ZN(n423) );
  NAND2_X1 U810 ( .A1(N155), .A2(n5750), .ZN(n425) );
  NAND2_X1 U811 ( .A1(N160), .A2(n5750), .ZN(n420) );
  NAND2_X1 U812 ( .A1(N162), .A2(n5760), .ZN(n418) );
  OAI21_X1 U813 ( .B1(n5800), .B2(n1450), .A(n416), .ZN(MB[19]) );
  NAND2_X1 U814 ( .A1(N164), .A2(n5760), .ZN(n416) );
  NAND2_X1 U815 ( .A1(N166), .A2(n5760), .ZN(n413) );
  OAI21_X1 U816 ( .B1(n579), .B2(n1550), .A(n403), .ZN(MB[9]) );
  NAND2_X1 U817 ( .A1(N154), .A2(n5750), .ZN(n403) );
  OAI21_X1 U818 ( .B1(n579), .B2(n1590), .A(n407), .ZN(MB[5]) );
  NAND2_X1 U819 ( .A1(N150), .A2(n5760), .ZN(n407) );
  NAND2_X1 U820 ( .A1(N148), .A2(n5760), .ZN(n409) );
  OAI21_X1 U821 ( .B1(n579), .B2(n1570), .A(n405), .ZN(MB[7]) );
  NAND2_X1 U822 ( .A1(N152), .A2(n5750), .ZN(n405) );
  OAI21_X1 U823 ( .B1(n5810), .B2(n1510), .A(n422), .ZN(MB[13]) );
  NAND2_X1 U824 ( .A1(N158), .A2(n5760), .ZN(n422) );
  OAI21_X1 U825 ( .B1(n5810), .B2(n1530), .A(n424), .ZN(MB[11]) );
  NAND2_X1 U826 ( .A1(N156), .A2(n5750), .ZN(n424) );
  OAI21_X1 U827 ( .B1(n5800), .B2(n1420), .A(n412), .ZN(MB[22]) );
  NAND2_X1 U828 ( .A1(N167), .A2(n5760), .ZN(n412) );
  INV_X1 U829 ( .A(n615), .ZN(n624) );
  OAI21_X1 U830 ( .B1(n5800), .B2(n1600), .A(n408), .ZN(MB[4]) );
  NAND2_X1 U831 ( .A1(N149), .A2(n577), .ZN(n408) );
  NAND2_X1 U832 ( .A1(N151), .A2(n5750), .ZN(n406) );
  OAI22_X1 U833 ( .A1(n579), .A2(n746), .B1(n5860), .B2(n1940), .ZN(MA[2]) );
  INV_X1 U834 ( .A(N179), .ZN(n746) );
  NAND2_X1 U835 ( .A1(n428), .A2(n429), .ZN(IBB) );
  NOR4_X1 U836 ( .A1(B_reg[30]), .A2(B_reg[29]), .A3(B_reg[28]), .A4(B_reg[27]), .ZN(n429) );
  NAND2_X1 U837 ( .A1(n430), .A2(n431), .ZN(IBA) );
  NOR4_X1 U838 ( .A1(A_reg[30]), .A2(A_reg[29]), .A3(A_reg[28]), .A4(A_reg[27]), .ZN(n431) );
  OAI21_X1 U839 ( .B1(n256), .B2(n764), .A(n257), .ZN(n441) );
  NAND2_X1 U840 ( .A1(overFlow), .A2(n5620), .ZN(n257) );
  NAND2_X1 U841 ( .A1(result[30]), .A2(n5620), .ZN(n336) );
  OAI21_X1 U842 ( .B1(n267), .B2(n764), .A(n341), .ZN(n437) );
  NAND2_X1 U843 ( .A1(result[25]), .A2(n5620), .ZN(n341) );
  OAI21_X1 U844 ( .B1(n266), .B2(n764), .A(n340), .ZN(n436) );
  NAND2_X1 U845 ( .A1(result[26]), .A2(n5620), .ZN(n340) );
  OAI21_X1 U846 ( .B1(n265), .B2(n764), .A(n339), .ZN(n435) );
  NAND2_X1 U847 ( .A1(result[27]), .A2(n5620), .ZN(n339) );
  OAI21_X1 U848 ( .B1(n264), .B2(n764), .A(n338), .ZN(n434) );
  NAND2_X1 U849 ( .A1(result[28]), .A2(n5620), .ZN(n338) );
  OAI21_X1 U850 ( .B1(n2010), .B2(n764), .A(n2020), .ZN(n439) );
  NAND2_X1 U851 ( .A1(result[23]), .A2(n5620), .ZN(n2020) );
  OAI21_X1 U852 ( .B1(n1980), .B2(n764), .A(n1990), .ZN(n438) );
  NAND2_X1 U853 ( .A1(result[24]), .A2(n5610), .ZN(n1990) );
  OAI21_X1 U854 ( .B1(n262), .B2(n764), .A(n337), .ZN(n433) );
  NAND2_X1 U855 ( .A1(result[29]), .A2(n5620), .ZN(n337) );
  OAI22_X1 U856 ( .A1(n579), .A2(n76), .B1(n588), .B2(n1660), .ZN(N208) );
  INV_X1 U857 ( .A(n345), .ZN(sub_78_B_2_) );
  INV_X1 U858 ( .A(n344), .ZN(sub_78_B_1_) );
  NAND2_X1 U859 ( .A1(N147), .A2(n5750), .ZN(n410) );
  INV_X1 U860 ( .A(n347), .ZN(sub_78_B_4_) );
  NAND2_X1 U861 ( .A1(n250), .A2(n251), .ZN(n440) );
  AOI22_X1 U862 ( .A1(N213), .A2(n522), .B1(result[0]), .B2(n5610), .ZN(n250)
         );
  AOI22_X1 U863 ( .A1(N549), .A2(n539), .B1(N212), .B2(n2050), .ZN(n251) );
  INV_X1 U864 ( .A(n334), .ZN(n738) );
  AOI22_X1 U865 ( .A1(n5620), .A2(result[31]), .B1(n335), .B2(enable), .ZN(
        n334) );
  OAI22_X1 U866 ( .A1(n74), .A2(n5630), .B1(n1650), .B2(n572), .ZN(n335) );
  OAI22_X1 U867 ( .A1(n578), .A2(n1390), .B1(n5830), .B2(n1710), .ZN(N203) );
  OAI22_X1 U868 ( .A1(n579), .A2(n1370), .B1(n5830), .B2(n1690), .ZN(N205) );
  OAI22_X1 U869 ( .A1(n578), .A2(n136), .B1(n5820), .B2(n1680), .ZN(N206) );
  INV_X1 U870 ( .A(enable), .ZN(n764) );
  NOR2_X1 U871 ( .A1(reset), .A2(enable), .ZN(n2000) );
  NAND2_X1 U872 ( .A1(A[23]), .A2(n548), .ZN(n2930) );
  NAND2_X1 U873 ( .A1(B[23]), .A2(n5510), .ZN(n3250) );
  NOR2_X1 U874 ( .A1(n764), .A2(reset), .ZN(n270) );
  OAI21_X1 U875 ( .B1(n1650), .B2(n5550), .A(n3010), .ZN(n473) );
  NAND2_X1 U876 ( .A1(A[31]), .A2(n5490), .ZN(n3010) );
  OAI21_X1 U877 ( .B1(n5580), .B2(n1960), .A(n269), .ZN(n442) );
  NAND2_X1 U878 ( .A1(A[0]), .A2(n547), .ZN(n269) );
  OAI21_X1 U879 ( .B1(n5570), .B2(n1950), .A(n271), .ZN(n443) );
  NAND2_X1 U880 ( .A1(A[1]), .A2(n547), .ZN(n271) );
  OAI21_X1 U881 ( .B1(n5570), .B2(n1920), .A(n274), .ZN(n446) );
  NAND2_X1 U882 ( .A1(A[4]), .A2(n547), .ZN(n274) );
  OAI21_X1 U883 ( .B1(n5570), .B2(n1890), .A(n277), .ZN(n449) );
  NAND2_X1 U884 ( .A1(A[7]), .A2(n547), .ZN(n277) );
  OAI21_X1 U885 ( .B1(n5570), .B2(n1870), .A(n279), .ZN(n451) );
  NAND2_X1 U886 ( .A1(A[9]), .A2(n547), .ZN(n279) );
  OAI21_X1 U887 ( .B1(n5570), .B2(n1860), .A(n2800), .ZN(n452) );
  NAND2_X1 U888 ( .A1(A[10]), .A2(n547), .ZN(n2800) );
  OAI21_X1 U889 ( .B1(n5570), .B2(n1850), .A(n2810), .ZN(n453) );
  NAND2_X1 U890 ( .A1(A[11]), .A2(n547), .ZN(n2810) );
  OAI21_X1 U891 ( .B1(n5570), .B2(n1840), .A(n2820), .ZN(n454) );
  NAND2_X1 U892 ( .A1(A[12]), .A2(n548), .ZN(n2820) );
  OAI21_X1 U893 ( .B1(n5580), .B2(n1830), .A(n2830), .ZN(n455) );
  NAND2_X1 U894 ( .A1(A[13]), .A2(n548), .ZN(n2830) );
  OAI21_X1 U895 ( .B1(n5570), .B2(n1820), .A(n2840), .ZN(n456) );
  NAND2_X1 U896 ( .A1(A[14]), .A2(n548), .ZN(n2840) );
  OAI21_X1 U897 ( .B1(n5580), .B2(n1810), .A(n2850), .ZN(n457) );
  NAND2_X1 U898 ( .A1(A[15]), .A2(n548), .ZN(n2850) );
  OAI21_X1 U899 ( .B1(n5570), .B2(n1800), .A(n2860), .ZN(n458) );
  NAND2_X1 U900 ( .A1(A[16]), .A2(n548), .ZN(n2860) );
  OAI21_X1 U901 ( .B1(n5570), .B2(n1790), .A(n2870), .ZN(n459) );
  NAND2_X1 U902 ( .A1(A[17]), .A2(n548), .ZN(n2870) );
  OAI21_X1 U903 ( .B1(n5570), .B2(n1780), .A(n2880), .ZN(n460) );
  NAND2_X1 U904 ( .A1(A[18]), .A2(n548), .ZN(n2880) );
  OAI21_X1 U905 ( .B1(n5580), .B2(n1770), .A(n2890), .ZN(n461) );
  NAND2_X1 U906 ( .A1(A[19]), .A2(n548), .ZN(n2890) );
  OAI21_X1 U907 ( .B1(n5570), .B2(n1760), .A(n2900), .ZN(n462) );
  NAND2_X1 U908 ( .A1(A[20]), .A2(n548), .ZN(n2900) );
  OAI21_X1 U909 ( .B1(n5570), .B2(n1750), .A(n2910), .ZN(n463) );
  NAND2_X1 U910 ( .A1(A[21]), .A2(n548), .ZN(n2910) );
  OAI21_X1 U911 ( .B1(n5580), .B2(n1740), .A(n2920), .ZN(n464) );
  NAND2_X1 U912 ( .A1(A[22]), .A2(n548), .ZN(n2920) );
  OAI21_X1 U913 ( .B1(n5580), .B2(n1640), .A(n3020), .ZN(n474) );
  NAND2_X1 U914 ( .A1(B[0]), .A2(n5490), .ZN(n3020) );
  OAI21_X1 U915 ( .B1(n5580), .B2(n1630), .A(n3030), .ZN(n475) );
  NAND2_X1 U916 ( .A1(B[1]), .A2(n5490), .ZN(n3030) );
  OAI21_X1 U917 ( .B1(n5580), .B2(n1620), .A(n3040), .ZN(n476) );
  NAND2_X1 U918 ( .A1(B[2]), .A2(n5490), .ZN(n3040) );
  OAI21_X1 U919 ( .B1(n5580), .B2(n1610), .A(n3050), .ZN(n477) );
  NAND2_X1 U920 ( .A1(B[3]), .A2(n5490), .ZN(n3050) );
  OAI21_X1 U921 ( .B1(n5580), .B2(n1600), .A(n3060), .ZN(n478) );
  NAND2_X1 U922 ( .A1(B[4]), .A2(n5500), .ZN(n3060) );
  OAI21_X1 U923 ( .B1(n5580), .B2(n1590), .A(n3070), .ZN(n479) );
  NAND2_X1 U924 ( .A1(B[5]), .A2(n5500), .ZN(n3070) );
  OAI21_X1 U925 ( .B1(n5580), .B2(n1580), .A(n3080), .ZN(n4800) );
  NAND2_X1 U926 ( .A1(B[6]), .A2(n5500), .ZN(n3080) );
  OAI21_X1 U927 ( .B1(n5580), .B2(n1570), .A(n3090), .ZN(n4810) );
  NAND2_X1 U928 ( .A1(B[7]), .A2(n5500), .ZN(n3090) );
  OAI21_X1 U929 ( .B1(n5590), .B2(n1560), .A(n3100), .ZN(n4820) );
  NAND2_X1 U930 ( .A1(B[8]), .A2(n5500), .ZN(n3100) );
  OAI21_X1 U931 ( .B1(n5590), .B2(n1550), .A(n3110), .ZN(n4830) );
  NAND2_X1 U932 ( .A1(B[9]), .A2(n5500), .ZN(n3110) );
  OAI21_X1 U933 ( .B1(n5590), .B2(n1540), .A(n3120), .ZN(n4840) );
  NAND2_X1 U934 ( .A1(B[10]), .A2(n5500), .ZN(n3120) );
  OAI21_X1 U935 ( .B1(n5590), .B2(n1530), .A(n3130), .ZN(n485) );
  NAND2_X1 U936 ( .A1(B[11]), .A2(n5500), .ZN(n3130) );
  OAI21_X1 U937 ( .B1(n5590), .B2(n1520), .A(n3140), .ZN(n486) );
  NAND2_X1 U938 ( .A1(B[12]), .A2(n5500), .ZN(n3140) );
  OAI21_X1 U939 ( .B1(n5590), .B2(n1510), .A(n3150), .ZN(n487) );
  NAND2_X1 U940 ( .A1(B[13]), .A2(n5500), .ZN(n3150) );
  OAI21_X1 U941 ( .B1(n5590), .B2(n1500), .A(n3160), .ZN(n488) );
  NAND2_X1 U942 ( .A1(B[14]), .A2(n5500), .ZN(n3160) );
  OAI21_X1 U943 ( .B1(n5590), .B2(n1490), .A(n3170), .ZN(n489) );
  NAND2_X1 U944 ( .A1(B[15]), .A2(n5500), .ZN(n3170) );
  OAI21_X1 U945 ( .B1(n5590), .B2(n1480), .A(n3180), .ZN(n490) );
  NAND2_X1 U946 ( .A1(B[16]), .A2(n5510), .ZN(n3180) );
  OAI21_X1 U947 ( .B1(n5590), .B2(n1470), .A(n3190), .ZN(n491) );
  NAND2_X1 U948 ( .A1(B[17]), .A2(n5510), .ZN(n3190) );
  OAI21_X1 U949 ( .B1(n5590), .B2(n1460), .A(n3200), .ZN(n492) );
  NAND2_X1 U950 ( .A1(B[18]), .A2(n5510), .ZN(n3200) );
  OAI21_X1 U951 ( .B1(n5590), .B2(n1450), .A(n3210), .ZN(n493) );
  NAND2_X1 U952 ( .A1(B[19]), .A2(n5510), .ZN(n3210) );
  OAI21_X1 U953 ( .B1(n5590), .B2(n1440), .A(n3220), .ZN(n494) );
  NAND2_X1 U954 ( .A1(B[20]), .A2(n5510), .ZN(n3220) );
  OAI21_X1 U955 ( .B1(n1400), .B2(n5550), .A(n3260), .ZN(n498) );
  NAND2_X1 U956 ( .A1(B[24]), .A2(n5510), .ZN(n3260) );
  OAI21_X1 U957 ( .B1(n1390), .B2(n5550), .A(n3270), .ZN(n499) );
  NAND2_X1 U958 ( .A1(B[25]), .A2(n5510), .ZN(n3270) );
  OAI21_X1 U959 ( .B1(n1380), .B2(n5550), .A(n328), .ZN(n500) );
  NAND2_X1 U960 ( .A1(B[26]), .A2(n5510), .ZN(n328) );
  OAI21_X1 U961 ( .B1(n1370), .B2(n5550), .A(n329), .ZN(n501) );
  NAND2_X1 U962 ( .A1(B[27]), .A2(n5510), .ZN(n329) );
  OAI21_X1 U963 ( .B1(n136), .B2(n5550), .A(n330), .ZN(n502) );
  NAND2_X1 U964 ( .A1(B[28]), .A2(n5520), .ZN(n330) );
  OAI21_X1 U965 ( .B1(n1350), .B2(n5550), .A(n331), .ZN(n503) );
  NAND2_X1 U966 ( .A1(B[29]), .A2(n5520), .ZN(n331) );
  OAI21_X1 U967 ( .B1(n76), .B2(n5550), .A(n332), .ZN(n504) );
  NAND2_X1 U968 ( .A1(B[30]), .A2(n5520), .ZN(n332) );
  OAI21_X1 U969 ( .B1(n1710), .B2(n5560), .A(n2950), .ZN(n467) );
  NAND2_X1 U970 ( .A1(A[25]), .A2(n5490), .ZN(n2950) );
  OAI21_X1 U971 ( .B1(n1700), .B2(n5560), .A(n2960), .ZN(n468) );
  NAND2_X1 U972 ( .A1(A[26]), .A2(n5490), .ZN(n2960) );
  OAI21_X1 U973 ( .B1(n1690), .B2(n5560), .A(n2970), .ZN(n469) );
  NAND2_X1 U974 ( .A1(A[27]), .A2(n5490), .ZN(n2970) );
  OAI21_X1 U975 ( .B1(n1680), .B2(n5560), .A(n2980), .ZN(n470) );
  NAND2_X1 U976 ( .A1(A[28]), .A2(n5490), .ZN(n2980) );
  OAI21_X1 U977 ( .B1(n1670), .B2(n5550), .A(n2990), .ZN(n471) );
  NAND2_X1 U978 ( .A1(A[29]), .A2(n5490), .ZN(n2990) );
  OAI21_X1 U979 ( .B1(n1660), .B2(n5560), .A(n3000), .ZN(n472) );
  NAND2_X1 U980 ( .A1(A[30]), .A2(n5490), .ZN(n3000) );
  OAI21_X1 U981 ( .B1(n1720), .B2(n5560), .A(n2940), .ZN(n466) );
  NAND2_X1 U982 ( .A1(A[24]), .A2(n5490), .ZN(n2940) );
  OAI21_X1 U983 ( .B1(n74), .B2(n5550), .A(n333), .ZN(n505) );
  NAND2_X1 U984 ( .A1(B[31]), .A2(n5520), .ZN(n333) );
  OAI21_X1 U985 ( .B1(n5560), .B2(n1940), .A(n272), .ZN(n444) );
  NAND2_X1 U986 ( .A1(A[2]), .A2(n547), .ZN(n272) );
  OAI21_X1 U987 ( .B1(n5560), .B2(n1930), .A(n273), .ZN(n445) );
  NAND2_X1 U988 ( .A1(A[3]), .A2(n547), .ZN(n273) );
  OAI21_X1 U989 ( .B1(n5560), .B2(n1910), .A(n275), .ZN(n447) );
  NAND2_X1 U990 ( .A1(A[5]), .A2(n547), .ZN(n275) );
  OAI21_X1 U991 ( .B1(n5560), .B2(n1900), .A(n276), .ZN(n448) );
  NAND2_X1 U992 ( .A1(A[6]), .A2(n547), .ZN(n276) );
  OAI21_X1 U993 ( .B1(n5560), .B2(n1880), .A(n2780), .ZN(n450) );
  NAND2_X1 U994 ( .A1(A[8]), .A2(n547), .ZN(n2780) );
  OAI21_X1 U995 ( .B1(n5560), .B2(n1420), .A(n3240), .ZN(n496) );
  NAND2_X1 U996 ( .A1(B[22]), .A2(n5510), .ZN(n3240) );
  OAI21_X1 U997 ( .B1(n5550), .B2(n1430), .A(n3230), .ZN(n495) );
  NAND2_X1 U998 ( .A1(B[21]), .A2(n5510), .ZN(n3230) );
  OR2_X1 U999 ( .A1(reset), .A2(n5520), .ZN(n268) );
  AOI22_X1 U1000 ( .A1(N215), .A2(n538), .B1(result[2]), .B2(n5610), .ZN(n247)
         );
  INV_X1 U1001 ( .A(n346), .ZN(n525) );
  INV_X1 U1002 ( .A(n346), .ZN(n526) );
  INV_X1 U1003 ( .A(n346), .ZN(N575) );
  INV_X1 U1004 ( .A(N575), .ZN(n605) );
  AOI21_X1 U1005 ( .B1(n342), .B2(MSB[0]), .A(N480), .ZN(n527) );
  OAI211_X1 U1006 ( .C1(n382), .C2(n383), .A(n381), .B(n520), .ZN(N481) );
  OAI21_X1 U1007 ( .B1(sll_78_A_22_), .B2(n393), .A(n520), .ZN(N480) );
  AOI22_X1 U1008 ( .A1(N327), .A2(n5640), .B1(N303), .B2(n5630), .ZN(n378) );
  OAI22_X1 U1009 ( .A1(n763), .A2(n577), .B1(n592), .B2(n1960), .ZN(MA[0]) );
  NOR2_X1 U1010 ( .A1(n516), .A2(n532), .ZN(n529) );
  CLKBUF_X1 U1011 ( .A(n261), .Z(n530) );
  INV_X1 U1012 ( .A(n528), .ZN(n672) );
  OAI22_X1 U1013 ( .A1(n579), .A2(n515), .B1(n5850), .B2(n1730), .ZN(N201) );
  AOI221_X1 U1014 ( .B1(n542), .B2(N559), .C1(n2050), .C2(N222), .A(n714), 
        .ZN(n2300) );
  INV_X1 U1015 ( .A(n1410), .ZN(n531) );
  OAI21_X1 U1016 ( .B1(n515), .B2(n5550), .A(n3250), .ZN(n497) );
  AOI221_X1 U1017 ( .B1(n540), .B2(N568), .C1(n2050), .C2(N231), .A(n732), 
        .ZN(n2120) );
  NOR2_X1 U1018 ( .A1(n255), .A2(n532), .ZN(n252) );
  NAND2_X1 U1019 ( .A1(enable), .A2(n765), .ZN(n532) );
  INV_X1 U1020 ( .A(n1730), .ZN(n533) );
  AOI221_X1 U1021 ( .B1(n539), .B2(N561), .C1(n543), .C2(N224), .A(n718), .ZN(
        n2260) );
  AOI221_X1 U1022 ( .B1(n540), .B2(N571), .C1(n2050), .C2(N234), .A(n737), 
        .ZN(n2030) );
  AOI221_X1 U1023 ( .B1(n542), .B2(N557), .C1(n543), .C2(N220), .A(n710), .ZN(
        n2340) );
  OAI21_X1 U1024 ( .B1(n1730), .B2(n5550), .A(n2930), .ZN(n465) );
  AOI221_X1 U1025 ( .B1(n541), .B2(N569), .C1(n544), .C2(N232), .A(n734), .ZN(
        n210) );
  AND2_X1 U1026 ( .A1(n253), .A2(n254), .ZN(n2040) );
  AND2_X1 U1027 ( .A1(n539), .A2(N570), .ZN(n534) );
  AND2_X1 U1028 ( .A1(n2050), .A2(N233), .ZN(n535) );
  BUF_X2 U1029 ( .A(n2040), .Z(n539) );
  INV_X1 U1030 ( .A(n209), .ZN(n735) );
  INV_X1 U1031 ( .A(n248), .ZN(n696) );
  INV_X1 U1032 ( .A(n2360), .ZN(n707) );
  INV_X1 U1033 ( .A(n2240), .ZN(n719) );
  AND2_X1 U1034 ( .A1(n542), .A2(N551), .ZN(n536) );
  AND2_X1 U1035 ( .A1(n2050), .A2(N214), .ZN(n537) );
  INV_X1 U1036 ( .A(n2450), .ZN(n700) );
  AOI221_X1 U1037 ( .B1(n541), .B2(N553), .C1(n544), .C2(N216), .A(n702), .ZN(
        n2420) );
  INV_X1 U1038 ( .A(n2430), .ZN(n702) );
  INV_X1 U1039 ( .A(n2310), .ZN(n714) );
  AOI221_X1 U1040 ( .B1(n540), .B2(N565), .C1(n543), .C2(N228), .A(n726), .ZN(
        n2180) );
  INV_X1 U1041 ( .A(n2190), .ZN(n726) );
  INV_X1 U1042 ( .A(n2130), .ZN(n732) );
  INV_X1 U1043 ( .A(n2320), .ZN(n711) );
  INV_X1 U1044 ( .A(n2200), .ZN(n723) );
  INV_X1 U1045 ( .A(n2400), .ZN(n703) );
  INV_X1 U1046 ( .A(n2280), .ZN(n715) );
  INV_X1 U1047 ( .A(n2160), .ZN(n727) );
  AOI221_X1 U1048 ( .B1(n540), .B2(N555), .C1(n544), .C2(N218), .A(n706), .ZN(
        n2380) );
  INV_X1 U1049 ( .A(n2390), .ZN(n706) );
  INV_X1 U1050 ( .A(n2270), .ZN(n718) );
  AOI221_X1 U1051 ( .B1(n542), .B2(N567), .C1(n543), .C2(N230), .A(n730), .ZN(
        n2140) );
  INV_X1 U1052 ( .A(n2150), .ZN(n730) );
  INV_X1 U1053 ( .A(n2350), .ZN(n710) );
  AOI221_X1 U1054 ( .B1(n540), .B2(N563), .C1(n543), .C2(N226), .A(n722), .ZN(
        n2220) );
  INV_X1 U1055 ( .A(n2230), .ZN(n722) );
  NOR2_X1 U1056 ( .A1(n258), .A2(n516), .ZN(n256) );
  INV_X1 U1057 ( .A(n211), .ZN(n734) );
  NOR2_X1 U1058 ( .A1(n764), .A2(n255), .ZN(n253) );
  AOI22_X1 U1059 ( .A1(n5210), .A2(N234), .B1(result[21]), .B2(n5600), .ZN(
        n209) );
  INV_X1 U1060 ( .A(n249), .ZN(n697) );
  AOI221_X1 U1061 ( .B1(n541), .B2(N550), .C1(n544), .C2(N213), .A(n697), .ZN(
        n248) );
  INV_X1 U1062 ( .A(n2420), .ZN(n701) );
  INV_X1 U1063 ( .A(n237), .ZN(n708) );
  AOI221_X1 U1064 ( .B1(n541), .B2(N556), .C1(n543), .C2(N219), .A(n708), .ZN(
        n2360) );
  INV_X1 U1065 ( .A(n2300), .ZN(n713) );
  INV_X1 U1066 ( .A(n2250), .ZN(n720) );
  AOI221_X1 U1067 ( .B1(n539), .B2(N562), .C1(n544), .C2(N225), .A(n720), .ZN(
        n2240) );
  AOI221_X1 U1068 ( .B1(n540), .B2(N552), .C1(n544), .C2(N215), .A(n700), .ZN(
        n2440) );
  AOI22_X1 U1069 ( .A1(N216), .A2(n5210), .B1(result[3]), .B2(n5610), .ZN(
        n2450) );
  INV_X1 U1070 ( .A(n2410), .ZN(n704) );
  AOI221_X1 U1071 ( .B1(n539), .B2(N554), .C1(n544), .C2(N217), .A(n704), .ZN(
        n2400) );
  INV_X1 U1072 ( .A(n2340), .ZN(n709) );
  INV_X1 U1073 ( .A(n2290), .ZN(n716) );
  AOI221_X1 U1074 ( .B1(n542), .B2(N560), .C1(n543), .C2(N223), .A(n716), .ZN(
        n2280) );
  INV_X1 U1075 ( .A(n2220), .ZN(n721) );
  INV_X1 U1076 ( .A(n2170), .ZN(n728) );
  AOI221_X1 U1077 ( .B1(n541), .B2(N566), .C1(n544), .C2(N229), .A(n728), .ZN(
        n2160) );
  INV_X1 U1078 ( .A(n2380), .ZN(n705) );
  INV_X1 U1079 ( .A(n2330), .ZN(n712) );
  AOI221_X1 U1080 ( .B1(n541), .B2(N558), .C1(n543), .C2(N221), .A(n712), .ZN(
        n2320) );
  INV_X1 U1081 ( .A(n2260), .ZN(n717) );
  INV_X1 U1082 ( .A(n2210), .ZN(n724) );
  AOI221_X1 U1083 ( .B1(n539), .B2(N564), .C1(n544), .C2(N227), .A(n724), .ZN(
        n2200) );
  INV_X1 U1084 ( .A(n2140), .ZN(n729) );
  INV_X1 U1085 ( .A(n2030), .ZN(n736) );
  INV_X1 U1086 ( .A(n2060), .ZN(n737) );
  NOR4_X1 U1087 ( .A1(B_reg[26]), .A2(B_reg[25]), .A3(B_reg[24]), .A4(n531), 
        .ZN(n428) );
  NAND2_X1 U1088 ( .A1(N145), .A2(n5750), .ZN(n426) );
  INV_X1 U1089 ( .A(n247), .ZN(n698) );
  NOR4_X1 U1090 ( .A1(A_reg[26]), .A2(A_reg[25]), .A3(A_reg[24]), .A4(n533), 
        .ZN(n430) );
  INV_X1 U1091 ( .A(n2440), .ZN(n699) );
  INV_X1 U1092 ( .A(n2180), .ZN(n725) );
  AOI22_X1 U1093 ( .A1(N232), .A2(n2070), .B1(result[19]), .B2(n5600), .ZN(
        n2130) );
  AOI22_X1 U1094 ( .A1(N229), .A2(n2070), .B1(result[16]), .B2(n5600), .ZN(
        n2190) );
  AOI22_X1 U1095 ( .A1(N226), .A2(n2070), .B1(result[13]), .B2(n5600), .ZN(
        n2250) );
  AOI22_X1 U1096 ( .A1(N223), .A2(n2070), .B1(result[10]), .B2(n5610), .ZN(
        n2310) );
  AOI22_X1 U1097 ( .A1(N220), .A2(n2070), .B1(result[7]), .B2(n5610), .ZN(n237) );
  AOI22_X1 U1098 ( .A1(N217), .A2(n2070), .B1(result[4]), .B2(n5610), .ZN(
        n2430) );
  AOI22_X1 U1099 ( .A1(N214), .A2(n2070), .B1(result[1]), .B2(n5610), .ZN(n249) );
  AND2_X1 U1100 ( .A1(n514), .A2(n351), .ZN(N483) );
  AND4_X2 U1101 ( .A1(n514), .A2(n348), .A3(n349), .A4(n350), .ZN(n342) );
  INV_X1 U1102 ( .A(n2120), .ZN(n731) );
  INV_X1 U1103 ( .A(n210), .ZN(n733) );
  AOI22_X1 U1104 ( .A1(N224), .A2(n538), .B1(result[11]), .B2(n5600), .ZN(
        n2290) );
  AOI22_X1 U1105 ( .A1(N233), .A2(n538), .B1(result[20]), .B2(n5600), .ZN(n211) );
  AOI22_X1 U1106 ( .A1(N230), .A2(n522), .B1(result[17]), .B2(n5600), .ZN(
        n2170) );
  AOI22_X1 U1107 ( .A1(N227), .A2(n5210), .B1(result[14]), .B2(n5600), .ZN(
        n2230) );
  AOI22_X1 U1108 ( .A1(N221), .A2(n538), .B1(result[8]), .B2(n5610), .ZN(n2350) );
  AOI22_X1 U1109 ( .A1(N218), .A2(n538), .B1(result[5]), .B2(n5610), .ZN(n2410) );
  NOR2_X1 U1110 ( .A1(n342), .A2(n765), .ZN(N612) );
  OAI21_X1 U1111 ( .B1(n530), .B2(n764), .A(n336), .ZN(n432) );
  AOI21_X1 U1112 ( .B1(n342), .B2(MSB[4]), .A(N484), .ZN(n347) );
  AOI21_X1 U1113 ( .B1(n342), .B2(MSB[2]), .A(N482), .ZN(n345) );
  AOI21_X1 U1114 ( .B1(n342), .B2(MSB[3]), .A(N483), .ZN(n346) );
  AOI21_X1 U1115 ( .B1(n342), .B2(MSB[1]), .A(N481), .ZN(n344) );
  INV_X1 U1116 ( .A(n358), .ZN(n739) );
  NOR2_X1 U1117 ( .A1(sll_78_A_16_), .A2(n358), .ZN(n357) );
  INV_X1 U1118 ( .A(N177), .ZN(n763) );
  AOI222_X1 U1119 ( .A1(N587), .A2(n254), .B1(n263), .B2(N208), .C1(N245), 
        .C2(n258), .ZN(n261) );
  AOI22_X1 U1120 ( .A1(N235), .A2(n538), .B1(result[22]), .B2(n5600), .ZN(
        n2060) );
  AOI22_X1 U1121 ( .A1(N231), .A2(n522), .B1(result[18]), .B2(n5600), .ZN(
        n2150) );
  AOI22_X1 U1122 ( .A1(N228), .A2(n5210), .B1(result[15]), .B2(n5600), .ZN(
        n2210) );
  AOI22_X1 U1123 ( .A1(N225), .A2(n538), .B1(result[12]), .B2(n5600), .ZN(
        n2270) );
  AOI22_X1 U1124 ( .A1(N222), .A2(n5210), .B1(result[9]), .B2(n5610), .ZN(
        n2330) );
  AOI22_X1 U1125 ( .A1(N219), .A2(n522), .B1(result[6]), .B2(n5610), .ZN(n2390) );
  AND2_X2 U1126 ( .A1(n252), .A2(N236), .ZN(n538) );
  BUF_X1 U1127 ( .A(n270), .Z(n545) );
  BUF_X1 U1128 ( .A(n270), .Z(n546) );
  BUF_X1 U1129 ( .A(n546), .Z(n5520) );
  BUF_X1 U1130 ( .A(n268), .Z(n5530) );
  BUF_X1 U1131 ( .A(n268), .Z(n5540) );
  BUF_X1 U1132 ( .A(N135), .Z(n574) );
  INV_X1 U1133 ( .A(n593), .ZN(n5810) );
  INV_X1 U1134 ( .A(n574), .ZN(n594) );
  INV_X1 U1135 ( .A(n574), .ZN(n595) );
  INV_X1 U1136 ( .A(n5810), .ZN(n596) );
  AND2_X1 U1137 ( .A1(sll_78_A_0_), .A2(n509), .ZN(sll_78_ML_int_1__0_) );
  AND2_X1 U1138 ( .A1(sll_78_ML_int_1__0_), .A2(sub_78_B_1_), .ZN(
        sll_78_ML_int_2__0_) );
  AND2_X1 U1139 ( .A1(sll_78_ML_int_1__1_), .A2(sub_78_B_1_), .ZN(
        sll_78_ML_int_2__1_) );
  AND2_X1 U1140 ( .A1(sll_78_ML_int_2__0_), .A2(sub_78_B_2_), .ZN(
        sll_78_ML_int_3__0_) );
  AND2_X1 U1141 ( .A1(sll_78_ML_int_2__1_), .A2(sub_78_B_2_), .ZN(
        sll_78_ML_int_3__1_) );
  AND2_X1 U1142 ( .A1(sll_78_ML_int_2__2_), .A2(sub_78_B_2_), .ZN(
        sll_78_ML_int_3__2_) );
  AND2_X1 U1143 ( .A1(sll_78_ML_int_2__3_), .A2(sub_78_B_2_), .ZN(
        sll_78_ML_int_3__3_) );
  NAND2_X1 U1144 ( .A1(sll_78_ML_int_3__0_), .A2(n605), .ZN(n597) );
  NAND2_X1 U1145 ( .A1(sll_78_ML_int_3__1_), .A2(n605), .ZN(n598) );
  NAND2_X1 U1146 ( .A1(sll_78_ML_int_3__2_), .A2(n605), .ZN(n599) );
  NAND2_X1 U1147 ( .A1(sll_78_ML_int_3__3_), .A2(n605), .ZN(n600) );
  NAND2_X1 U1148 ( .A1(sll_78_ML_int_3__4_), .A2(n605), .ZN(n601) );
  NAND2_X1 U1149 ( .A1(sll_78_ML_int_3__5_), .A2(n605), .ZN(n602) );
  NAND2_X1 U1150 ( .A1(sll_78_ML_int_3__6_), .A2(n605), .ZN(n603) );
  NAND2_X1 U1151 ( .A1(n606), .A2(n508), .ZN(n604) );
  NOR2_X1 U1152 ( .A1(n604), .A2(n597), .ZN(N549) );
  AND2_X1 U1153 ( .A1(sll_78_ML_int_4__10_), .A2(n607), .ZN(N559) );
  AND2_X1 U1154 ( .A1(sll_78_ML_int_4__11_), .A2(n607), .ZN(N560) );
  AND2_X1 U1155 ( .A1(sll_78_ML_int_4__12_), .A2(n607), .ZN(N561) );
  AND2_X1 U1156 ( .A1(sll_78_ML_int_4__13_), .A2(n607), .ZN(N562) );
  AND2_X1 U1157 ( .A1(sll_78_ML_int_4__14_), .A2(n607), .ZN(N563) );
  AND2_X1 U1158 ( .A1(sll_78_ML_int_4__15_), .A2(n607), .ZN(N564) );
  AND2_X1 U1159 ( .A1(sll_78_ML_int_5__16_), .A2(n508), .ZN(N565) );
  AND2_X1 U1160 ( .A1(sll_78_ML_int_5__17_), .A2(n508), .ZN(N566) );
  AND2_X1 U1161 ( .A1(sll_78_ML_int_5__18_), .A2(n508), .ZN(N567) );
  AND2_X1 U1162 ( .A1(sll_78_ML_int_5__19_), .A2(n508), .ZN(N568) );
  NOR2_X1 U1163 ( .A1(n604), .A2(n598), .ZN(N550) );
  AND2_X1 U1164 ( .A1(sll_78_ML_int_5__20_), .A2(n508), .ZN(N569) );
  AND2_X1 U1165 ( .A1(sll_78_ML_int_5__21_), .A2(n508), .ZN(N570) );
  AND2_X1 U1166 ( .A1(sll_78_ML_int_5__22_), .A2(n508), .ZN(N571) );
  NOR2_X1 U1167 ( .A1(n604), .A2(n599), .ZN(N551) );
  NOR2_X1 U1168 ( .A1(n604), .A2(n600), .ZN(N552) );
  NOR2_X1 U1169 ( .A1(n604), .A2(n601), .ZN(N553) );
  NOR2_X1 U1170 ( .A1(n604), .A2(n602), .ZN(N554) );
  NOR2_X1 U1171 ( .A1(n604), .A2(n603), .ZN(N555) );
  AND3_X1 U1172 ( .A1(n607), .A2(n605), .A3(sll_78_ML_int_3__7_), .ZN(N556) );
  AND2_X1 U1173 ( .A1(sll_78_ML_int_4__8_), .A2(n607), .ZN(N557) );
  AND2_X1 U1174 ( .A1(sll_78_ML_int_4__9_), .A2(n607), .ZN(N558) );
  NOR2_X1 U1175 ( .A1(B_reg[29]), .A2(n1670), .ZN(n622) );
  NOR2_X1 U1176 ( .A1(n1730), .A2(n531), .ZN(n615) );
  AOI21_X1 U1177 ( .B1(n615), .B2(n1400), .A(A_reg[24]), .ZN(n616) );
  AOI221_X1 U1178 ( .B1(B_reg[25]), .B2(n1710), .C1(B_reg[24]), .C2(n624), .A(
        n616), .ZN(n617) );
  AOI221_X1 U1179 ( .B1(A_reg[26]), .B2(n1380), .C1(A_reg[25]), .C2(n1390), 
        .A(n617), .ZN(n618) );
  AOI221_X1 U1180 ( .B1(B_reg[27]), .B2(n1690), .C1(B_reg[26]), .C2(n1700), 
        .A(n618), .ZN(n619) );
  AOI221_X1 U1181 ( .B1(A_reg[28]), .B2(n136), .C1(A_reg[27]), .C2(n1370), .A(
        n619), .ZN(n620) );
  AOI221_X1 U1182 ( .B1(B_reg[29]), .B2(n1670), .C1(B_reg[28]), .C2(n1680), 
        .A(n620), .ZN(n621) );
  OAI22_X1 U1183 ( .A1(n622), .A2(n621), .B1(A_reg[30]), .B2(n76), .ZN(n623)
         );
  OAI21_X1 U1184 ( .B1(B_reg[30]), .B2(n1660), .A(n623), .ZN(N135) );
  OAI211_X1 U1185 ( .C1(MB[1]), .C2(n687), .A(n672), .B(n5180), .ZN(n625) );
  OAI221_X1 U1186 ( .B1(MA[1]), .B2(n665), .C1(MA[2]), .C2(n666), .A(n625), 
        .ZN(n626) );
  OAI221_X1 U1187 ( .B1(MB[2]), .B2(n688), .C1(MB[3]), .C2(n689), .A(n626), 
        .ZN(n627) );
  OAI221_X1 U1188 ( .B1(MA[3]), .B2(n667), .C1(MA[4]), .C2(n671), .A(n627), 
        .ZN(n628) );
  OAI221_X1 U1189 ( .B1(MB[4]), .B2(n693), .C1(MB[5]), .C2(n692), .A(n628), 
        .ZN(n629) );
  OAI221_X1 U1190 ( .B1(MA[5]), .B2(n670), .C1(MA[6]), .C2(n669), .A(n629), 
        .ZN(n630) );
  OAI221_X1 U1191 ( .B1(MB[6]), .B2(n691), .C1(MB[7]), .C2(n690), .A(n630), 
        .ZN(n631) );
  OAI221_X1 U1192 ( .B1(MA[7]), .B2(n668), .C1(MA[8]), .C2(n654), .A(n631), 
        .ZN(n632) );
  OAI221_X1 U1193 ( .B1(MB[8]), .B2(n678), .C1(MB[9]), .C2(n677), .A(n632), 
        .ZN(n633) );
  OAI221_X1 U1194 ( .B1(MA[10]), .B2(n664), .C1(MA[9]), .C2(n653), .A(n633), 
        .ZN(n634) );
  OAI221_X1 U1195 ( .B1(MB[10]), .B2(n686), .C1(MB[11]), .C2(n685), .A(n634), 
        .ZN(n635) );
  OAI221_X1 U1196 ( .B1(MA[11]), .B2(n663), .C1(MA[12]), .C2(n662), .A(n635), 
        .ZN(n636) );
  OAI221_X1 U1197 ( .B1(MB[12]), .B2(n684), .C1(MB[13]), .C2(n683), .A(n636), 
        .ZN(n637) );
  OAI221_X1 U1198 ( .B1(MA[13]), .B2(n661), .C1(MA[14]), .C2(n660), .A(n637), 
        .ZN(n638) );
  OAI221_X1 U1199 ( .B1(MB[14]), .B2(n682), .C1(MB[15]), .C2(n681), .A(n638), 
        .ZN(n639) );
  OAI221_X1 U1200 ( .B1(MA[15]), .B2(n659), .C1(MA[16]), .C2(n652), .A(n639), 
        .ZN(n640) );
  OAI221_X1 U1201 ( .B1(MB[16]), .B2(n676), .C1(MB[17]), .C2(n675), .A(n640), 
        .ZN(n641) );
  OAI221_X1 U1202 ( .B1(MA[17]), .B2(n651), .C1(MA[18]), .C2(n650), .A(n641), 
        .ZN(n642) );
  OAI221_X1 U1203 ( .B1(MB[18]), .B2(n674), .C1(MB[19]), .C2(n673), .A(n642), 
        .ZN(n643) );
  OAI221_X1 U1204 ( .B1(MA[19]), .B2(n649), .C1(MA[20]), .C2(n658), .A(n643), 
        .ZN(n644) );
  OAI221_X1 U1205 ( .B1(MB[20]), .B2(n680), .C1(MB[21]), .C2(n679), .A(n644), 
        .ZN(n645) );
  OAI221_X1 U1206 ( .B1(MA[21]), .B2(n657), .C1(MA[22]), .C2(n656), .A(n645), 
        .ZN(n646) );
  AOI21_X1 U1207 ( .B1(n656), .B2(MA[22]), .A(n694), .ZN(n648) );
  OAI21_X1 U1208 ( .B1(n695), .B2(n655), .A(r145_B_23_), .ZN(n647) );
  OAI21_X1 U1209 ( .B1(MB[23]), .B2(n648), .A(n647), .ZN(N278) );
endmodule

